magic
tech sky130A
timestamp 1702422646
<< nwell >>
rect -125 20 945 1770
<< pmos >>
rect 0 905 50 1505
rect 100 905 150 1505
rect 285 905 335 1505
rect 485 905 535 1505
rect 670 905 720 1505
rect 770 905 820 1505
rect 0 75 50 675
rect 100 75 150 675
rect 200 75 250 675
rect 570 75 620 675
rect 670 75 720 675
rect 770 75 820 675
<< pdiff >>
rect -50 1490 0 1505
rect -50 920 -35 1490
rect -15 920 0 1490
rect -50 905 0 920
rect 50 1490 100 1505
rect 50 920 65 1490
rect 85 920 100 1490
rect 50 905 100 920
rect 150 1490 200 1505
rect 150 920 165 1490
rect 185 920 200 1490
rect 150 905 200 920
rect 235 1490 285 1505
rect 235 920 250 1490
rect 270 920 285 1490
rect 235 905 285 920
rect 335 1490 385 1505
rect 335 920 350 1490
rect 370 920 385 1490
rect 335 905 385 920
rect 435 1490 485 1505
rect 435 920 450 1490
rect 470 920 485 1490
rect 435 905 485 920
rect 535 1490 585 1505
rect 535 920 550 1490
rect 570 920 585 1490
rect 535 905 585 920
rect 620 1490 670 1505
rect 620 920 635 1490
rect 655 920 670 1490
rect 620 905 670 920
rect 720 1490 770 1505
rect 720 920 735 1490
rect 755 920 770 1490
rect 720 905 770 920
rect 820 1490 870 1505
rect 820 920 835 1490
rect 855 920 870 1490
rect 820 905 870 920
rect -50 660 0 675
rect -50 90 -35 660
rect -15 90 0 660
rect -50 75 0 90
rect 50 660 100 675
rect 50 90 65 660
rect 85 90 100 660
rect 50 75 100 90
rect 150 660 200 675
rect 150 90 165 660
rect 185 90 200 660
rect 150 75 200 90
rect 250 660 300 675
rect 250 90 265 660
rect 285 90 300 660
rect 520 660 570 675
rect 250 75 300 90
rect 520 90 535 660
rect 555 90 570 660
rect 520 75 570 90
rect 620 660 670 675
rect 620 90 635 660
rect 655 90 670 660
rect 620 75 670 90
rect 720 660 770 675
rect 720 90 735 660
rect 755 90 770 660
rect 720 75 770 90
rect 820 660 870 675
rect 820 90 835 660
rect 855 90 870 660
rect 820 75 870 90
<< pdiffc >>
rect -35 920 -15 1490
rect 65 920 85 1490
rect 165 920 185 1490
rect 250 920 270 1490
rect 350 920 370 1490
rect 450 920 470 1490
rect 550 920 570 1490
rect 635 920 655 1490
rect 735 920 755 1490
rect 835 920 855 1490
rect -35 90 -15 660
rect 65 90 85 660
rect 165 90 185 660
rect 265 90 285 660
rect 535 90 555 660
rect 635 90 655 660
rect 735 90 755 660
rect 835 90 855 660
<< nsubdiff >>
rect -100 1495 -50 1505
rect -100 920 -85 1495
rect -65 920 -50 1495
rect -100 905 -50 920
rect 870 1495 920 1505
rect 870 920 885 1495
rect 905 920 920 1495
rect 870 905 920 920
rect -100 665 -50 675
rect -100 90 -85 665
rect -65 90 -50 665
rect -100 75 -50 90
rect 870 665 920 675
rect 870 90 885 665
rect 905 90 920 665
rect 870 75 920 90
<< nsubdiffcont >>
rect -85 920 -65 1495
rect 885 920 905 1495
rect -85 90 -65 665
rect 885 90 905 665
<< poly >>
rect 190 1700 240 1710
rect 190 1680 200 1700
rect 220 1680 240 1700
rect 190 1675 240 1680
rect 580 1700 630 1710
rect 580 1680 600 1700
rect 620 1680 630 1700
rect 580 1675 630 1680
rect 50 1650 80 1660
rect 50 1630 55 1650
rect 75 1640 80 1650
rect 140 1650 170 1660
rect 140 1640 145 1650
rect 75 1630 145 1640
rect 165 1630 170 1650
rect 50 1625 170 1630
rect 50 1620 80 1625
rect 140 1620 170 1625
rect 100 1550 150 1560
rect 100 1530 110 1550
rect 130 1530 150 1550
rect 0 1505 50 1520
rect 100 1505 150 1530
rect 0 890 50 905
rect 100 890 150 905
rect 0 880 35 890
rect 0 860 5 880
rect 25 860 35 880
rect 210 860 225 1675
rect 285 1650 335 1660
rect 285 1630 295 1650
rect 315 1630 335 1650
rect 285 1625 335 1630
rect 485 1650 535 1660
rect 485 1630 505 1650
rect 525 1630 535 1650
rect 485 1625 535 1630
rect 285 1520 300 1625
rect 520 1520 535 1625
rect 285 1505 335 1520
rect 485 1505 535 1520
rect 285 890 335 905
rect 485 890 535 905
rect 0 850 35 860
rect 135 845 225 860
rect 595 860 610 1675
rect 650 1650 680 1660
rect 650 1630 655 1650
rect 675 1640 680 1650
rect 740 1650 770 1660
rect 740 1640 745 1650
rect 675 1630 745 1640
rect 765 1630 770 1650
rect 650 1625 770 1630
rect 650 1620 680 1625
rect 740 1620 770 1625
rect 670 1550 720 1560
rect 670 1530 690 1550
rect 710 1530 720 1550
rect 670 1505 720 1530
rect 770 1505 820 1520
rect 670 890 720 905
rect 770 890 820 905
rect 785 880 820 890
rect 785 860 795 880
rect 815 860 820 880
rect 595 845 685 860
rect 785 850 820 860
rect 100 840 150 845
rect 100 820 110 840
rect 130 820 150 840
rect 100 810 150 820
rect 670 840 720 845
rect 670 820 690 840
rect 710 820 720 840
rect 670 810 720 820
rect -30 780 20 790
rect -30 760 -20 780
rect 0 770 20 780
rect 800 780 850 790
rect 800 770 820 780
rect 0 760 820 770
rect 840 760 850 780
rect -30 755 850 760
rect 100 720 150 730
rect 100 700 110 720
rect 130 700 150 720
rect 0 675 50 690
rect 100 675 150 700
rect 200 690 215 755
rect 380 720 430 730
rect 380 700 390 720
rect 410 700 430 720
rect 380 695 430 700
rect 200 675 250 690
rect 400 630 415 695
rect 605 690 620 755
rect 570 675 620 690
rect 670 720 720 730
rect 670 700 690 720
rect 710 700 720 720
rect 670 675 720 700
rect 770 675 820 690
rect 380 620 430 630
rect 380 600 390 620
rect 410 600 430 620
rect 380 595 430 600
rect 0 60 50 75
rect 100 60 150 75
rect 200 60 250 75
rect 570 60 620 75
rect 670 60 720 75
rect 770 60 820 75
rect 0 50 35 60
rect 0 30 5 50
rect 25 30 35 50
rect 0 20 35 30
rect 785 50 820 60
rect 785 30 795 50
rect 815 30 820 50
rect 785 20 820 30
<< polycont >>
rect 200 1680 220 1700
rect 600 1680 620 1700
rect 55 1630 75 1650
rect 145 1630 165 1650
rect 110 1530 130 1550
rect 5 860 25 880
rect 295 1630 315 1650
rect 505 1630 525 1650
rect 655 1630 675 1650
rect 745 1630 765 1650
rect 690 1530 710 1550
rect 795 860 815 880
rect 110 820 130 840
rect 690 820 710 840
rect -20 760 0 780
rect 820 760 840 780
rect 110 700 130 720
rect 390 700 410 720
rect 690 700 710 720
rect 390 600 410 620
rect 5 30 25 50
rect 795 30 815 50
<< locali >>
rect 50 1650 80 1660
rect 50 1645 55 1650
rect -125 1630 55 1645
rect 75 1630 80 1650
rect -125 1625 80 1630
rect 50 1620 80 1625
rect 100 1600 120 1770
rect 205 1750 225 1770
rect 205 1730 615 1750
rect 205 1710 225 1730
rect 595 1710 615 1730
rect 190 1700 240 1710
rect 190 1680 200 1700
rect 220 1680 240 1700
rect 190 1675 240 1680
rect 580 1700 630 1710
rect 580 1680 600 1700
rect 620 1680 630 1700
rect 580 1675 630 1680
rect 140 1650 170 1660
rect 140 1630 145 1650
rect 165 1645 170 1650
rect 285 1650 335 1660
rect 285 1645 295 1650
rect 165 1630 295 1645
rect 315 1645 335 1650
rect 485 1650 535 1660
rect 485 1645 505 1650
rect 315 1630 505 1645
rect 525 1645 535 1650
rect 650 1650 680 1660
rect 650 1645 655 1650
rect 525 1630 655 1645
rect 675 1630 680 1650
rect 140 1625 680 1630
rect 140 1620 170 1625
rect 650 1620 680 1625
rect 740 1650 770 1660
rect 740 1630 745 1650
rect 765 1645 770 1650
rect 765 1630 945 1645
rect 740 1625 945 1630
rect 740 1620 770 1625
rect 100 1580 720 1600
rect 100 1560 120 1580
rect 700 1560 720 1580
rect 100 1550 150 1560
rect 100 1530 110 1550
rect 130 1530 150 1550
rect 100 1520 150 1530
rect 670 1550 720 1560
rect 670 1530 690 1550
rect 710 1530 720 1550
rect 670 1520 720 1530
rect -95 1495 -5 1500
rect -95 920 -85 1495
rect -65 920 -35 1495
rect -15 920 -5 1495
rect -95 910 -5 920
rect -25 890 -5 910
rect 55 1490 95 1500
rect 55 920 65 1490
rect 85 920 95 1490
rect 55 910 95 920
rect 155 1495 195 1500
rect 155 920 165 1495
rect 185 920 195 1495
rect 155 910 195 920
rect 240 1490 280 1500
rect 240 920 250 1490
rect 270 920 280 1490
rect 240 910 280 920
rect 340 1490 380 1500
rect 340 920 350 1490
rect 370 930 380 1490
rect 440 1490 480 1500
rect 440 930 450 1490
rect 370 920 450 930
rect 470 920 480 1490
rect 340 910 480 920
rect 540 1490 580 1500
rect 540 920 550 1490
rect 570 920 580 1490
rect 540 910 580 920
rect 625 1495 665 1500
rect 625 920 635 1495
rect 655 920 665 1495
rect 625 910 665 920
rect 725 1490 765 1500
rect 725 920 735 1490
rect 755 920 765 1490
rect 725 910 765 920
rect -25 880 35 890
rect -25 870 5 880
rect 0 860 5 870
rect 25 860 35 880
rect 0 850 35 860
rect -30 780 20 790
rect -30 775 -20 780
rect -125 760 -20 775
rect 0 760 20 780
rect -125 755 20 760
rect 55 670 75 910
rect 240 890 260 910
rect 175 870 260 890
rect 100 840 150 845
rect 100 820 110 840
rect 130 820 150 840
rect 100 810 150 820
rect 130 730 150 810
rect 100 720 150 730
rect 100 700 110 720
rect 130 700 150 720
rect 100 690 150 700
rect 175 670 195 870
rect 400 730 420 910
rect 560 890 580 910
rect 560 870 645 890
rect 380 720 430 730
rect 380 700 390 720
rect 410 700 430 720
rect 380 695 430 700
rect 625 670 645 870
rect 670 840 720 845
rect 670 820 690 840
rect 710 820 720 840
rect 670 810 720 820
rect 670 730 690 810
rect 670 720 720 730
rect 670 700 690 720
rect 710 700 720 720
rect 670 690 720 700
rect 745 670 765 910
rect 825 1495 915 1500
rect 825 920 835 1495
rect 855 920 885 1495
rect 905 920 915 1495
rect 825 910 915 920
rect 825 890 845 910
rect 785 880 845 890
rect 785 860 795 880
rect 815 870 845 880
rect 815 860 820 870
rect 785 850 820 860
rect 800 780 850 790
rect 800 760 820 780
rect 840 775 850 780
rect 840 760 945 775
rect 800 755 945 760
rect -95 665 -5 670
rect -95 90 -85 665
rect -65 90 -35 665
rect -15 90 -5 665
rect -95 80 -5 90
rect 55 660 95 670
rect 55 90 65 660
rect 85 90 95 660
rect 55 80 95 90
rect 155 660 195 670
rect 155 90 165 660
rect 185 90 195 660
rect 155 80 195 90
rect 255 660 565 670
rect 255 90 265 660
rect 285 650 535 660
rect 285 90 295 650
rect 255 80 295 90
rect -25 60 -5 80
rect -25 50 35 60
rect -25 40 5 50
rect 0 30 5 40
rect 25 30 35 50
rect 0 20 35 30
rect 320 20 340 650
rect 380 620 430 630
rect 380 600 390 620
rect 410 600 430 620
rect 380 595 430 600
rect 390 20 410 595
rect 525 90 535 650
rect 555 90 565 660
rect 525 80 565 90
rect 625 660 665 670
rect 625 90 635 660
rect 655 90 665 660
rect 625 80 665 90
rect 725 660 765 670
rect 725 90 735 660
rect 755 90 765 660
rect 725 80 765 90
rect 825 665 915 670
rect 825 90 835 665
rect 855 90 885 665
rect 905 90 915 665
rect 825 80 915 90
rect 825 60 845 80
rect 785 50 845 60
rect 785 30 795 50
rect 815 40 845 50
rect 815 30 820 40
rect 785 20 820 30
<< viali >>
rect -85 920 -65 1495
rect -35 1490 -15 1495
rect -35 920 -15 1490
rect 165 1490 185 1495
rect 165 920 185 1490
rect 635 1490 655 1495
rect 635 920 655 1490
rect 835 1490 855 1495
rect 835 920 855 1490
rect 885 920 905 1495
rect -85 90 -65 665
rect -35 660 -15 665
rect -35 90 -15 660
rect 835 660 855 665
rect 835 90 855 660
rect 885 90 905 665
<< metal1 >>
rect -125 1495 945 1500
rect -125 920 -85 1495
rect -65 920 -35 1495
rect -15 920 165 1495
rect 185 920 635 1495
rect 655 920 835 1495
rect 855 920 885 1495
rect 905 920 945 1495
rect -125 665 945 920
rect -125 90 -85 665
rect -65 90 -35 665
rect -15 90 835 665
rect 855 90 885 665
rect 905 90 945 665
rect -125 80 945 90
<< labels >>
rlabel locali -125 765 -125 765 7 Vphi
port 1 w
rlabel locali -125 1635 -125 1635 7 Vphi_b
port 2 w
rlabel locali 110 1770 110 1770 1 Vbp
port 3 n
rlabel locali 215 1770 215 1770 1 Vcp
port 4 n
rlabel locali 330 20 330 20 5 Viun
port 5 s
rlabel locali 400 20 400 20 5 Viup
port 6 s
rlabel metal1 -125 1495 -125 1495 7 VP
port 7 w
<< end >>
