* NGSPICE file created from final.ext - technology: sky130A

.subckt v_gen VP VN Vb Vcp Vbp
X0 VP VP Vcp VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X1 VP VP Vbp VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X2 VN Vb a_500_1500# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X3 a_800_1390# a_800_1390# a_2400_1500# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X4 a_800_1390# a_800_1390# a_2400_1500# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X5 VN VN Vbp VN sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X6 a_2640_60# Vb a_2440_60# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X7 VN Vb a_2840_60# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X8 VN Vb Vb VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X9 VN Vb Vbp VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X10 a_2240_60# Vb a_800_1390# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X11 VP Vbp Vbp VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X12 a_800_1390# Vb a_1660_60# VN sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X13 a_700_1500# a_500_1500# a_500_1500# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X14 a_700_1500# a_800_1390# a_800_1390# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X15 a_1460_60# Vb a_1260_60# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X16 a_700_1500# a_800_1390# a_800_1390# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X17 Vbp VN VN VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X18 Vcp Vcp a_2400_1500# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X19 Vbp Vbp VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X20 a_1060_60# Vb VN VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X21 a_2400_1500# a_800_1390# VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X22 a_2400_1500# a_800_1390# a_800_1390# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X23 Vb Vb VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X24 a_2840_60# Vb a_2640_60# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X25 Vbp Vb VN VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X26 a_2440_60# Vb a_2240_60# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X27 Vbp VP VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X28 a_500_1500# VP VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X29 a_1660_60# Vb a_1460_60# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X30 a_800_1390# a_800_1390# a_700_1500# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X31 a_800_1390# a_800_1390# a_700_1500# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X32 a_1260_60# Vb a_1060_60# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X33 VP a_800_1390# a_700_1500# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X34 a_2400_1500# a_800_1390# a_800_1390# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X35 Vcp Vb VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
.ends

.subckt dac_unit Vphi Vphi_b Vbp Vcp Viun Viup VP
X0 a_1440_150# Vcp a_1070_1810# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X1 VP Vbp a_100_150# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X2 a_1440_150# Vbp VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X3 a_300_150# Vcp a_100_150# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X4 Viup Vphi_b a_300_150# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=3 ps=13 w=6 l=0.5
X5 a_1070_1810# Vphi_b Viup VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=3 ps=13 w=6 l=0.5
X6 VP VP a_1440_150# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X7 a_100_150# VP VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X8 a_1070_1810# Vphi Viun VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X9 a_100_150# VP VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X10 Viun Vphi a_300_150# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X11 VP VP a_1440_150# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
.ends

.subckt inverter A Y VP VN
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
.ends

.subckt dac_v2 Vcp Vphi1 Vphi2 Vphi3 Vphi4 Vphi5 Vphi6 Vphi7 Viout- Viout+ Vbp inverter_7/VP
+ VSUBS
Xdac_unit_4 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_5 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_6 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xinverter_0 Vphi7 inverter_0/Y inverter_7/VP VSUBS inverter
Xinverter_1 Vphi2 inverter_1/Y inverter_7/VP VSUBS inverter
Xdac_unit_7 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_8 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xinverter_2 Vphi3 inverter_2/Y inverter_7/VP VSUBS inverter
Xinverter_3 Vphi4 inverter_3/Y inverter_7/VP VSUBS inverter
Xdac_unit_9 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xinverter_4 Vphi5 inverter_4/Y inverter_7/VP VSUBS inverter
Xinverter_5 Vphi6 inverter_5/Y inverter_7/VP VSUBS inverter
Xinverter_7 Vphi1 inverter_7/Y inverter_7/VP VSUBS inverter
Xdac_unit_40 Vphi1 inverter_7/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_41 Vphi1 inverter_7/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_30 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_42 Vphi1 inverter_7/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_20 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_31 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_10 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_21 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_32 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_11 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_22 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_33 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_12 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_23 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_34 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_14 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_13 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_25 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_24 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_36 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_35 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_15 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_26 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_16 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_27 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_17 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_28 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_18 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_29 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_19 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_0 Vphi7 inverter_0/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_1 Vphi7 inverter_0/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_3 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_2 Vphi7 inverter_0/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
.ends

.subckt filter VN Viout- Viout+
X0 Viout+ a_2360_6260# VN sky130_fd_pr__res_xhigh_po l=3.5
X1 VN a_2360_6260# VN sky130_fd_pr__res_xhigh_po l=3.5
X2 VN a_2360_1100# VN sky130_fd_pr__res_xhigh_po l=3.5
X3 a_1460_5820# a_1090_2450# sky130_fd_pr__cap_mim_m3_1 l=10 w=8
X4 Viout- a_2360_1100# VN sky130_fd_pr__res_xhigh_po l=3.5
X5 a_1460_5820# Vout+ VN sky130_fd_pr__res_xhigh_po l=3.5
X6 a_1090_2450# Viout- VN sky130_fd_pr__res_xhigh_po l=3.5
X7 a_1090_2450# Vout- VN sky130_fd_pr__res_xhigh_po l=3.5
X8 a_1460_5820# Viout+ VN sky130_fd_pr__res_xhigh_po l=3.5
X9 Vout+ Vout- sky130_fd_pr__cap_mim_m3_1 l=10 w=8
.ends

.subckt csrl_dff2 D DB Q QB CLK VP VN
X0 VP a_n950_630# a_n950_1180# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X1 a_n950_630# a_n950_1180# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X2 a_n950_630# CLK DB VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.75 ps=3.5 w=1 l=0.15
X3 QB CLK a_n950_630# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 VP a_n950_1180# a_n950_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X5 VN Q QB VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X6 a_n690_630# CLK VP VP sky130_fd_pr__pfet_01v8 ad=0.433 pd=3.03 as=0.5 ps=3.16 w=4 l=0.15
X7 a_n950_n280# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0.433 pd=3.03 as=2 ps=10.5 w=4 l=0.15
X8 a_n950_1180# a_n950_630# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X9 Q CLK a_n950_1180# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 VN QB Q VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X11 Q QB a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X12 QB Q a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X13 a_n950_1180# CLK D VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.75 ps=3.5 w=1 l=0.15
.ends

.subckt csrl_dff3 D DB Q QB CLK VP VN
X0 VP a_n950_630# a_n950_1180# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X1 a_n950_630# a_n950_1180# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X2 a_n950_630# CLK DB VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.75 ps=3.5 w=1 l=0.15
X3 QB CLK a_n950_630# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 VP a_n950_1180# a_n950_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X5 VN Q QB VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X6 a_n690_630# CLK VP VP sky130_fd_pr__pfet_01v8 ad=0.433 pd=3.03 as=0.5 ps=3.16 w=4 l=0.15
X7 a_n950_n280# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0.433 pd=3.03 as=2 ps=10.5 w=4 l=0.15
X8 a_n950_1180# a_n950_630# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X9 Q CLK a_n950_1180# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 VN QB Q VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X11 Q QB a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X12 QB Q a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X13 a_n950_1180# CLK D VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.75 ps=3.5 w=1 l=0.15
.ends

.subckt csrl_dff1 D DB Q QB CLK VP VN
X0 VP a_n950_630# a_n950_1180# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X1 a_n950_630# a_n950_1180# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X2 a_n950_630# CLK DB VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.55 ps=3.1 w=1 l=0.15
X3 QB CLK a_n950_630# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 VP a_n950_1180# a_n950_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X5 VN Q QB VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X6 a_n690_630# CLK VP VP sky130_fd_pr__pfet_01v8 ad=0.433 pd=3.03 as=0.5 ps=3.16 w=4 l=0.15
X7 a_n950_n280# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0.433 pd=3.03 as=1.6 ps=9.7 w=4 l=0.15
X8 a_n950_1180# a_n950_630# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X9 Q CLK a_n950_1180# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 VN QB Q VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X11 Q QB a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X12 QB Q a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X13 a_n950_1180# CLK D VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.55 ps=3.1 w=1 l=0.15
.ends

.subckt register16 Vphi3 csrl_dff3_0/VP Vphi7 Vphi1 Vphi5 Vphi2 Vphi4 Vphi6 VSUBS
Xcsrl_dff2_10 csrl_dff2_9/Q csrl_dff2_9/QB csrl_dff2_11/D csrl_dff2_11/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_11 csrl_dff2_11/D csrl_dff2_11/DB csrl_dff2_12/D csrl_dff2_12/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_12 csrl_dff2_12/D csrl_dff2_12/DB csrl_dff2_13/D csrl_dff2_13/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_0 Vphi1 csrl_dff2_0/DB Vphi2 csrl_dff2_1/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_13 csrl_dff2_13/D csrl_dff2_13/DB csrl_dff3_0/D csrl_dff3_0/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_2 Vphi3 csrl_dff2_2/DB Vphi4 csrl_dff2_3/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_1 Vphi2 csrl_dff2_1/DB Vphi3 csrl_dff2_2/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_3 Vphi4 csrl_dff2_3/DB Vphi5 csrl_dff2_4/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_4 Vphi5 csrl_dff2_4/DB Vphi6 csrl_dff2_5/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_5 Vphi6 csrl_dff2_5/DB Vphi7 csrl_dff2_6/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_6 Vphi7 csrl_dff2_6/DB csrl_dff2_7/D csrl_dff2_7/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_7 csrl_dff2_7/D csrl_dff2_7/DB csrl_dff2_8/D csrl_dff2_8/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_8 csrl_dff2_8/D csrl_dff2_8/DB csrl_dff2_9/D csrl_dff2_9/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_9 csrl_dff2_9/D csrl_dff2_9/DB csrl_dff2_9/Q csrl_dff2_9/QB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff3_0 csrl_dff3_0/D csrl_dff3_0/DB csrl_dff3_0/Q csrl_dff3_0/QB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff3
Xcsrl_dff1_0 csrl_dff3_0/Q csrl_dff3_0/QB Vphi1 csrl_dff2_0/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff1
.ends


* Top level circuit final

Xv_gen_0 v_gen_0/VP VSUBS v_gen_0/Vb v_gen_0/Vcp v_gen_0/Vbp v_gen
Xdac_v2_0 v_gen_0/Vcp dac_v2_0/Vphi1 dac_v2_0/Vphi2 dac_v2_0/Vphi3 dac_v2_0/Vphi4
+ dac_v2_0/Vphi5 dac_v2_0/Vphi6 dac_v2_0/Vphi7 filter_0/Viout- filter_0/Viout+ v_gen_0/Vbp
+ v_gen_0/VP VSUBS dac_v2
Xfilter_0 VSUBS filter_0/Viout- filter_0/Viout+ filter
Xregister16_0 dac_v2_0/Vphi3 v_gen_0/VP dac_v2_0/Vphi7 dac_v2_0/Vphi1 dac_v2_0/Vphi5
+ dac_v2_0/Vphi2 dac_v2_0/Vphi4 dac_v2_0/Vphi6 VSUBS register16
.end

