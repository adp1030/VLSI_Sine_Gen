magic
tech sky130A
timestamp 1702679324
<< nwell >>
rect -565 295 -220 805
<< nmos >>
rect -490 -140 -475 260
rect -435 160 -420 260
rect -370 160 -355 260
rect -305 160 -290 260
rect -435 -115 -420 -15
rect -370 -115 -355 -15
rect -305 -115 -290 -15
<< pmos >>
rect -490 590 -475 690
rect -425 590 -410 690
rect -490 315 -475 415
rect -425 315 -410 415
rect -360 315 -345 715
rect -305 590 -290 690
rect -305 315 -290 415
<< ndiff >>
rect -545 245 -490 260
rect -545 175 -530 245
rect -510 175 -490 245
rect -545 160 -490 175
rect -515 -15 -490 160
rect -545 -30 -490 -15
rect -545 -100 -530 -30
rect -510 -100 -490 -30
rect -545 -115 -490 -100
rect -515 -140 -490 -115
rect -475 160 -435 260
rect -420 245 -370 260
rect -420 175 -405 245
rect -385 175 -370 245
rect -420 160 -370 175
rect -355 245 -305 260
rect -355 175 -340 245
rect -320 175 -305 245
rect -355 160 -305 175
rect -290 245 -240 260
rect -290 175 -275 245
rect -255 175 -240 245
rect -290 160 -240 175
rect -475 -15 -450 160
rect -475 -115 -435 -15
rect -420 -30 -370 -15
rect -420 -100 -405 -30
rect -385 -100 -370 -30
rect -420 -115 -370 -100
rect -355 -30 -305 -15
rect -355 -100 -340 -30
rect -320 -100 -305 -30
rect -355 -115 -305 -100
rect -290 -30 -240 -15
rect -290 -100 -275 -30
rect -255 -100 -240 -30
rect -290 -115 -240 -100
rect -475 -140 -450 -115
<< pdiff >>
rect -385 690 -360 715
rect -545 675 -490 690
rect -545 605 -530 675
rect -510 605 -490 675
rect -545 590 -490 605
rect -475 675 -425 690
rect -475 605 -460 675
rect -440 605 -425 675
rect -475 590 -425 605
rect -410 675 -360 690
rect -410 605 -395 675
rect -375 605 -360 675
rect -410 590 -360 605
rect -385 415 -360 590
rect -545 400 -490 415
rect -545 330 -530 400
rect -510 330 -490 400
rect -545 315 -490 330
rect -475 400 -425 415
rect -475 330 -460 400
rect -440 330 -425 400
rect -475 315 -425 330
rect -410 400 -360 415
rect -410 330 -395 400
rect -375 330 -360 400
rect -410 315 -360 330
rect -345 690 -320 715
rect -345 590 -305 690
rect -290 675 -240 690
rect -290 605 -275 675
rect -255 605 -240 675
rect -290 590 -240 605
rect -345 415 -320 590
rect -345 315 -305 415
rect -290 400 -240 415
rect -290 330 -275 400
rect -255 330 -240 400
rect -290 315 -240 330
<< ndiffc >>
rect -530 175 -510 245
rect -530 -100 -510 -30
rect -405 175 -385 245
rect -340 175 -320 245
rect -275 175 -255 245
rect -405 -100 -385 -30
rect -340 -100 -320 -30
rect -275 -100 -255 -30
<< pdiffc >>
rect -530 605 -510 675
rect -460 605 -440 675
rect -395 605 -375 675
rect -530 330 -510 400
rect -460 330 -440 400
rect -395 330 -375 400
rect -275 605 -255 675
rect -275 330 -255 400
<< psubdiff >>
rect -370 -180 -255 -165
rect -370 -200 -350 -180
rect -275 -200 -255 -180
rect -370 -215 -255 -200
<< nsubdiff >>
rect -520 770 -405 785
rect -520 750 -500 770
rect -425 750 -405 770
rect -520 735 -405 750
<< psubdiffcont >>
rect -350 -200 -275 -180
<< nsubdiffcont >>
rect -500 750 -425 770
<< poly >>
rect -360 715 -345 730
rect -490 690 -475 705
rect -425 690 -410 705
rect -490 415 -475 590
rect -425 575 -410 590
rect -440 565 -400 575
rect -440 545 -430 565
rect -410 545 -400 565
rect -440 535 -400 545
rect -450 500 -410 510
rect -450 480 -440 500
rect -420 480 -410 500
rect -450 470 -410 480
rect -425 415 -410 470
rect -305 690 -290 705
rect -305 545 -290 590
rect -305 535 -265 545
rect -305 515 -295 535
rect -275 515 -265 535
rect -305 505 -265 515
rect -285 465 -245 475
rect -285 450 -275 465
rect -305 445 -275 450
rect -255 445 -245 465
rect -305 435 -245 445
rect -305 415 -290 435
rect -490 260 -475 315
rect -425 285 -410 315
rect -360 285 -345 315
rect -435 270 -410 285
rect -370 270 -345 285
rect -435 260 -420 270
rect -370 260 -355 270
rect -305 260 -290 315
rect -435 145 -420 160
rect -370 145 -355 160
rect -440 135 -400 145
rect -440 115 -430 135
rect -410 115 -400 135
rect -440 105 -400 115
rect -375 130 -355 145
rect -305 145 -290 160
rect -305 135 -255 145
rect -305 130 -285 135
rect -440 70 -400 80
rect -440 50 -430 70
rect -410 50 -400 70
rect -440 40 -400 50
rect -435 -15 -420 40
rect -375 10 -360 130
rect -295 115 -285 130
rect -265 115 -255 135
rect -295 105 -255 115
rect -335 70 -295 80
rect -335 50 -325 70
rect -305 50 -295 70
rect -335 40 -295 50
rect -310 10 -295 40
rect -375 -5 -355 10
rect -310 -5 -290 10
rect -370 -15 -355 -5
rect -305 -15 -290 -5
rect -435 -130 -420 -115
rect -370 -125 -355 -115
rect -395 -140 -355 -125
rect -305 -130 -290 -115
rect -490 -245 -475 -140
rect -395 -245 -380 -140
rect -490 -255 -450 -245
rect -490 -275 -480 -255
rect -460 -275 -450 -255
rect -490 -285 -450 -275
rect -420 -255 -380 -245
rect -420 -275 -410 -255
rect -390 -275 -380 -255
rect -420 -285 -380 -275
<< polycont >>
rect -430 545 -410 565
rect -440 480 -420 500
rect -295 515 -275 535
rect -275 445 -255 465
rect -430 115 -410 135
rect -430 50 -410 70
rect -285 115 -265 135
rect -325 50 -305 70
rect -480 -275 -460 -255
rect -410 -275 -390 -255
<< locali >>
rect -515 770 -410 780
rect -515 750 -500 770
rect -425 765 -410 770
rect -425 750 -385 765
rect -515 740 -385 750
rect -410 735 -385 740
rect -405 685 -385 735
rect -285 685 -265 805
rect -540 675 -500 685
rect -540 615 -530 675
rect -565 605 -530 615
rect -510 605 -500 675
rect -470 675 -430 685
rect -470 615 -460 675
rect -565 595 -500 605
rect -480 605 -460 615
rect -440 605 -430 675
rect -480 595 -430 605
rect -405 675 -365 685
rect -405 605 -395 675
rect -375 605 -365 675
rect -405 595 -365 605
rect -285 675 -245 685
rect -285 605 -275 675
rect -255 615 -245 675
rect -255 605 -225 615
rect -285 595 -225 605
rect -480 510 -460 595
rect -440 565 -400 575
rect -440 545 -430 565
rect -410 555 -400 565
rect -410 545 -370 555
rect -440 535 -370 545
rect -480 500 -410 510
rect -480 490 -440 500
rect -450 480 -440 490
rect -420 480 -410 500
rect -450 470 -410 480
rect -390 450 -370 535
rect -305 535 -265 545
rect -305 530 -295 535
rect -450 430 -370 450
rect -330 515 -295 530
rect -275 515 -265 535
rect -330 505 -265 515
rect -450 410 -430 430
rect -330 410 -310 505
rect -245 475 -225 595
rect -285 465 -225 475
rect -285 445 -275 465
rect -255 455 -225 465
rect -255 445 -245 455
rect -285 435 -245 445
rect -540 400 -500 410
rect -540 340 -530 400
rect -565 330 -530 340
rect -510 330 -500 400
rect -565 320 -500 330
rect -470 400 -430 410
rect -470 330 -460 400
rect -440 330 -430 400
rect -470 320 -430 330
rect -405 400 -365 410
rect -405 330 -395 400
rect -375 330 -365 400
rect -405 320 -365 330
rect -330 400 -245 410
rect -330 390 -275 400
rect -460 255 -440 320
rect -330 255 -310 390
rect -285 330 -275 390
rect -255 330 -245 400
rect -285 320 -245 330
rect -540 245 -500 255
rect -540 175 -530 245
rect -510 175 -500 245
rect -540 165 -500 175
rect -480 245 -375 255
rect -480 235 -405 245
rect -480 80 -460 235
rect -415 175 -405 235
rect -385 175 -375 245
rect -415 165 -375 175
rect -350 245 -310 255
rect -350 175 -340 245
rect -320 175 -310 245
rect -350 165 -310 175
rect -285 245 -245 255
rect -285 175 -275 245
rect -255 175 -245 245
rect -285 165 -245 175
rect -440 135 -400 145
rect -440 115 -430 135
rect -410 125 -400 135
rect -410 115 -360 125
rect -440 105 -360 115
rect -480 70 -400 80
rect -480 60 -430 70
rect -440 50 -430 60
rect -410 50 -400 70
rect -440 40 -400 50
rect -380 10 -360 105
rect -335 80 -315 165
rect -295 135 -255 145
rect -295 115 -285 135
rect -265 115 -255 135
rect -295 105 -255 115
rect -335 70 -295 80
rect -335 50 -325 70
rect -305 50 -295 70
rect -335 40 -295 50
rect -275 20 -255 105
rect -395 -5 -360 10
rect -330 0 -255 20
rect -395 -20 -370 -5
rect -330 -20 -310 0
rect -540 -30 -500 -20
rect -540 -100 -530 -30
rect -510 -100 -500 -30
rect -540 -110 -500 -100
rect -415 -30 -370 -20
rect -350 -30 -310 -20
rect -415 -100 -405 -30
rect -385 -100 -375 -30
rect -415 -110 -375 -100
rect -350 -100 -340 -30
rect -320 -100 -310 -30
rect -350 -110 -310 -100
rect -285 -30 -245 -20
rect -285 -100 -275 -30
rect -255 -100 -245 -30
rect -285 -110 -245 -100
rect -285 -170 -265 -110
rect -365 -180 -260 -170
rect -365 -200 -350 -180
rect -275 -200 -260 -180
rect -365 -210 -260 -200
rect -490 -255 -450 -245
rect -490 -275 -480 -255
rect -460 -275 -450 -255
rect -490 -285 -450 -275
rect -420 -255 -380 -245
rect -420 -275 -410 -255
rect -390 -275 -380 -255
rect -420 -285 -380 -275
<< viali >>
rect -500 750 -425 770
rect -395 605 -375 675
rect -395 330 -375 400
rect -530 175 -510 245
rect -275 175 -255 245
rect -530 -100 -510 -30
rect -275 -100 -255 -30
rect -350 -200 -275 -180
rect -480 -275 -460 -255
rect -410 -275 -390 -255
<< metal1 >>
rect -545 770 -240 785
rect -545 750 -500 770
rect -425 750 -240 770
rect -545 675 -240 750
rect -545 605 -395 675
rect -375 605 -240 675
rect -545 400 -240 605
rect -545 330 -395 400
rect -375 330 -240 400
rect -545 315 -240 330
rect -545 245 -240 260
rect -545 175 -530 245
rect -510 175 -275 245
rect -255 175 -240 245
rect -545 -30 -240 175
rect -545 -100 -530 -30
rect -510 -100 -275 -30
rect -255 -100 -240 -30
rect -545 -180 -240 -100
rect -545 -200 -350 -180
rect -275 -200 -240 -180
rect -370 -215 -255 -200
rect -545 -255 -240 -245
rect -545 -275 -480 -255
rect -460 -275 -410 -255
rect -390 -275 -240 -255
rect -545 -285 -240 -275
<< labels >>
rlabel metal1 -545 550 -545 550 7 VP
port 6 w
rlabel metal1 -545 45 -545 45 7 VN
port 7 w
rlabel locali -565 605 -565 605 7 D
port 1 w
rlabel locali -565 330 -565 330 7 DB
port 2 w
rlabel locali -275 805 -275 805 1 Q
port 3 n
rlabel locali -245 365 -245 365 3 QB
port 4 e
rlabel metal1 -545 -265 -545 -265 1 CLK
port 5 n
<< end >>
