magic
tech sky130A
timestamp 1702883810
<< psubdiff >>
rect 1385 1830 1535 1845
rect 1385 1800 1400 1830
rect 1520 1800 1535 1830
rect 1385 1785 1535 1800
rect 1530 1035 1590 1050
rect 1530 915 1545 1035
rect 1575 915 1590 1035
rect 1530 900 1590 915
rect 710 630 770 645
rect -250 595 -190 610
rect -250 475 -235 595
rect -205 475 -190 595
rect 710 510 725 630
rect 755 510 770 630
rect 710 495 770 510
rect -250 460 -190 475
<< psubdiffcont >>
rect 1400 1800 1520 1830
rect 1545 915 1575 1035
rect -235 475 -205 595
rect 725 510 755 630
<< xpolycontact >>
rect 715 1700 935 1735
rect 1285 1700 1505 1735
rect 1640 1225 1675 1445
rect -375 795 -155 830
rect 195 795 415 830
rect -375 690 -155 725
rect 195 690 415 725
rect 1640 655 1675 875
rect -135 575 85 610
rect 435 575 655 610
rect -135 515 85 550
rect 435 515 655 550
rect 820 610 1040 645
rect 1390 610 1610 645
rect 820 550 1040 585
rect 1390 550 1610 585
<< xpolyres >>
rect 935 1700 1285 1735
rect 1640 875 1675 1225
rect -155 795 195 830
rect -155 690 195 725
rect 85 575 435 610
rect 85 515 435 550
rect 1040 610 1390 645
rect 1040 550 1390 585
<< locali >>
rect 550 1735 590 1890
rect 1390 1830 1530 1840
rect 1390 1800 1400 1830
rect 1520 1800 1530 1830
rect 1390 1790 1530 1800
rect 445 1700 715 1735
rect 1505 1700 1675 1735
rect 445 1410 490 1700
rect 1640 1655 1675 1700
rect 540 1640 620 1655
rect 540 1540 555 1640
rect 605 1540 620 1640
rect 540 1525 620 1540
rect 1595 1640 1675 1655
rect 1595 1540 1610 1640
rect 1660 1540 1675 1640
rect 1595 1525 1675 1540
rect 1640 1445 1675 1525
rect 445 1395 570 1410
rect 445 1295 505 1395
rect 555 1295 570 1395
rect 445 1280 570 1295
rect 1535 1035 1585 1045
rect 490 1000 570 1015
rect 490 900 505 1000
rect 555 900 570 1000
rect 1535 915 1545 1035
rect 1575 915 1585 1035
rect 1535 905 1585 915
rect 490 890 570 900
rect -420 855 570 890
rect 195 830 570 855
rect 415 795 570 830
rect -375 780 -155 795
rect -375 750 -360 780
rect -240 750 -155 780
rect -375 725 -155 750
rect 415 690 655 725
rect 195 655 655 690
rect -420 630 655 655
rect 1640 645 1675 655
rect 435 610 655 630
rect -245 595 -195 605
rect -245 475 -235 595
rect -205 475 -195 595
rect 715 630 765 640
rect -135 550 85 575
rect -245 465 -195 475
rect 435 500 585 515
rect 715 510 725 630
rect 755 510 765 630
rect 1610 610 1685 645
rect 820 585 1040 610
rect 715 500 765 510
rect 1390 535 1540 550
rect 1390 505 1405 535
rect 1525 505 1540 535
rect 435 470 450 500
rect 570 470 585 500
rect 1390 490 1540 505
rect 435 455 585 470
<< viali >>
rect 1400 1800 1520 1830
rect 555 1540 605 1640
rect 1610 1540 1660 1640
rect 505 1295 555 1395
rect 505 900 555 1000
rect 1545 915 1575 1035
rect -360 750 -240 780
rect -235 475 -205 595
rect 725 510 755 630
rect 1405 505 1525 535
rect 450 470 570 500
<< metal1 >>
rect 1305 1830 1570 1865
rect 1305 1800 1400 1830
rect 1520 1800 1570 1830
rect 1305 1780 1570 1800
rect 540 1640 620 1655
rect 540 1540 555 1640
rect 605 1540 620 1640
rect 540 1525 620 1540
rect 1530 1475 1570 1780
rect 1595 1640 1675 1655
rect 1595 1540 1610 1640
rect 1660 1540 1675 1640
rect 1595 1525 1675 1540
rect 490 1395 570 1410
rect 490 1295 505 1395
rect 555 1295 570 1395
rect 490 1280 570 1295
rect 1530 1035 1590 1475
rect 490 1000 570 1015
rect 490 900 505 1000
rect 555 900 570 1000
rect 490 885 570 900
rect 1530 915 1545 1035
rect 1575 915 1590 1035
rect -375 780 -225 795
rect -375 750 -360 780
rect -240 750 -225 780
rect -375 735 -225 750
rect 1530 650 1590 915
rect -370 635 1590 650
rect -370 630 1595 635
rect -370 595 725 630
rect -370 475 -235 595
rect -205 510 725 595
rect 755 535 1595 630
rect 755 510 1405 535
rect -205 505 1405 510
rect 1525 505 1595 535
rect -205 500 1595 505
rect -205 475 450 500
rect -370 470 450 475
rect 570 470 1595 500
rect -370 455 1595 470
<< via1 >>
rect 555 1540 605 1640
rect 1610 1540 1660 1640
rect 505 1295 555 1395
rect 505 900 555 1000
rect -360 750 -240 780
<< metal2 >>
rect 540 1640 675 1655
rect 540 1540 555 1640
rect 605 1540 675 1640
rect 540 1525 675 1540
rect 1595 1640 1675 1655
rect 1595 1540 1610 1640
rect 1660 1540 1675 1640
rect 1595 1525 1675 1540
rect 490 1395 570 1410
rect 490 1295 505 1395
rect 555 1295 570 1395
rect 490 1280 570 1295
rect 490 1000 570 1015
rect 490 900 505 1000
rect 555 900 570 1000
rect 490 885 570 900
rect 600 795 675 1525
rect -375 780 675 795
rect -375 750 -360 780
rect -240 750 675 780
rect -375 735 675 750
<< via2 >>
rect 555 1540 605 1640
rect 1610 1540 1660 1640
rect 505 1295 555 1395
rect 505 900 555 1000
<< metal3 >>
rect -415 1410 425 1890
rect 690 1655 1520 1685
rect 540 1640 620 1655
rect 540 1540 555 1640
rect 605 1540 620 1640
rect 540 1525 620 1540
rect 690 1640 1675 1655
rect 690 1540 1610 1640
rect 1660 1540 1675 1640
rect 690 1525 1675 1540
rect -415 1395 570 1410
rect -415 1295 505 1395
rect 555 1295 570 1395
rect -415 1280 570 1295
rect -415 850 425 1280
rect 490 1000 570 1015
rect 490 900 505 1000
rect 555 900 570 1000
rect 490 885 570 900
rect 690 655 1520 1525
<< via3 >>
rect 555 1540 605 1640
rect 505 900 555 1000
<< mimcap >>
rect -395 1000 405 1870
rect -395 900 295 1000
rect 375 900 405 1000
rect -395 870 405 900
rect 705 1640 1505 1670
rect 705 1540 735 1640
rect 815 1540 1505 1640
rect 705 670 1505 1540
<< mimcapcontact >>
rect 295 900 375 1000
rect 735 1540 815 1640
<< metal4 >>
rect 540 1640 830 1655
rect 540 1540 555 1640
rect 605 1540 735 1640
rect 815 1540 830 1640
rect 540 1525 830 1540
rect 280 1000 570 1015
rect 280 900 295 1000
rect 375 900 505 1000
rect 555 900 570 1000
rect 280 885 570 900
<< labels >>
rlabel locali 1685 625 1685 625 3 Viout-
rlabel locali -420 640 -420 640 7 Viout+
rlabel locali 570 1890 570 1890 1 Vout-
rlabel locali -420 870 -420 870 7 Vout+
rlabel metal1 1305 1820 1305 1820 7 VN
<< end >>
