magic
tech sky130A
timestamp 1702440739
<< poly >>
rect -205 880 -165 890
rect -205 860 -195 880
rect -175 860 -165 880
rect -205 850 -165 860
rect 5325 880 5365 890
rect 5325 860 5335 880
rect 5355 860 5365 880
rect 5325 850 5365 860
rect -210 580 -170 590
rect -210 560 -200 580
rect -180 560 -170 580
rect -210 550 -170 560
rect 5330 580 5370 590
rect 5330 560 5340 580
rect 5360 560 5370 580
rect 5330 550 5370 560
<< polycont >>
rect -195 860 -175 880
rect 5335 860 5355 880
rect -200 560 -180 580
rect 5340 560 5360 580
<< locali >>
rect -205 880 -165 890
rect -205 860 -195 880
rect -175 870 -165 880
rect 5325 880 5365 890
rect 5325 870 5335 880
rect -175 860 -115 870
rect -205 850 -115 860
rect 175 850 225 870
rect 515 850 565 870
rect 855 850 905 870
rect 1195 850 1245 870
rect 1535 850 1585 870
rect 1875 850 1925 870
rect 2215 850 2265 870
rect 2555 850 2605 870
rect 2895 850 2945 870
rect 3235 850 3285 870
rect 3575 850 3625 870
rect 3915 850 3965 870
rect 4255 850 4305 870
rect 4595 850 4645 870
rect 4935 850 4985 870
rect 5275 860 5335 870
rect 5355 860 5365 880
rect 5275 850 5365 860
rect -210 580 -170 590
rect -210 560 -200 580
rect -180 570 -170 580
rect 5330 580 5370 590
rect 5330 570 5340 580
rect -180 560 -115 570
rect -210 550 -115 560
rect 175 550 225 570
rect 515 550 565 570
rect 855 550 905 570
rect 1195 550 1245 570
rect 1535 550 1585 570
rect 1875 550 1925 570
rect 2215 550 2265 570
rect 2555 550 2605 570
rect 2895 550 2945 570
rect 3235 550 3285 570
rect 3575 550 3625 570
rect 3915 550 3965 570
rect 4255 550 4305 570
rect 4595 550 4645 570
rect 4935 550 4985 570
rect 5275 560 5340 570
rect 5360 560 5370 580
rect 5275 550 5370 560
<< viali >>
rect -195 860 -175 880
rect 5335 860 5355 880
rect -200 560 -180 580
rect 5340 560 5360 580
<< metal1 >>
rect -235 1095 -220 1205
rect -235 1080 5395 1095
rect -235 585 -220 1080
rect -200 1050 5360 1065
rect -200 880 -170 1050
rect -200 860 -195 880
rect -175 860 -170 880
rect -200 850 -170 860
rect -265 580 -170 585
rect -265 560 -200 580
rect -180 560 -170 580
rect -265 555 -170 560
rect -140 545 -120 1020
rect 200 545 220 1020
rect 540 545 560 1020
rect 880 545 900 1020
rect 1220 545 1240 1020
rect 1560 545 1580 1020
rect 1900 545 1920 1020
rect 2240 545 2260 1020
rect 2580 545 2600 1020
rect 2920 545 2940 1020
rect 3260 545 3280 1020
rect 3600 545 3620 1020
rect 3940 545 3960 1020
rect 4280 545 4300 1020
rect 4620 545 4640 1020
rect 4960 545 4980 1020
rect 5330 880 5360 1050
rect 5330 860 5335 880
rect 5355 860 5360 880
rect 5330 850 5360 860
rect 5380 585 5395 1080
rect 5330 580 5395 585
rect 5330 560 5340 580
rect 5360 560 5395 580
rect 5330 555 5395 560
rect -140 40 -120 490
rect 200 40 220 490
rect 540 40 560 490
rect 880 40 900 490
rect 1220 40 1240 490
rect 1560 40 1580 490
rect 1900 40 1920 490
rect 2240 40 2260 490
rect 2580 40 2600 490
rect 2920 40 2940 490
rect 3260 40 3280 490
rect 3600 40 3620 490
rect 3940 40 3960 490
rect 4280 40 4300 490
rect 4620 40 4640 490
rect 4960 40 4980 490
rect -140 -30 -120 10
rect 200 -30 220 10
rect 540 -30 560 10
rect 880 -30 900 10
rect 1220 -30 1240 10
rect 1560 -30 1580 10
rect 1900 -30 1920 10
rect 2240 -30 2260 10
rect 2580 -30 2600 10
rect 2920 -30 2940 10
rect 3260 -30 3280 10
rect 3600 -30 3620 10
rect 3940 -30 3960 10
rect 4280 -30 4300 10
rect 4620 -30 4640 10
rect 4960 -30 4980 10
use csrl_dff  csrl_dff_0 ~/VLSI_Sine_Gen/layout/shift_register
timestamp 1695756208
transform 1 0 -90 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_2
timestamp 1695756208
transform 1 0 590 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_3
timestamp 1695756208
transform 1 0 930 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_4
timestamp 1695756208
transform 1 0 1270 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_5
timestamp 1695756208
transform 1 0 1610 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_6
timestamp 1695756208
transform 1 0 1950 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_7
timestamp 1695756208
transform 1 0 2290 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_8
timestamp 1695756208
transform 1 0 2630 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_9
timestamp 1695756208
transform 1 0 2970 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_10
timestamp 1695756208
transform 1 0 3310 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_11
timestamp 1695756208
transform 1 0 3650 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_12
timestamp 1695756208
transform 1 0 3990 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_13
timestamp 1695756208
transform 1 0 4330 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_14
timestamp 1695756208
transform 1 0 4670 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_15
timestamp 1695756208
transform 1 0 5010 0 1 230
box -50 -260 290 810
use csrl_dff  csrl_dff_16
timestamp 1695756208
transform 1 0 250 0 1 230
box -50 -260 290 810
<< end >>
