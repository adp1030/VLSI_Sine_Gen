magic
tech sky130A
timestamp 1702708471
<< metal3 >>
rect 700 3155 1530 3185
rect 625 3025 1530 3155
rect 700 2155 1530 3025
rect 700 1655 1530 1685
rect 625 1525 1530 1655
rect 700 655 1530 1525
<< mimcap >>
rect 715 3140 1515 3170
rect 715 3040 1405 3140
rect 1485 3040 1515 3140
rect 715 2170 1515 3040
rect 715 1640 1515 1670
rect 715 1540 1405 1640
rect 1485 1540 1515 1640
rect 715 670 1515 1540
<< mimcapcontact >>
rect 1405 3040 1485 3140
rect 1405 1540 1485 1640
<< metal4 >>
rect 1390 3140 1600 3155
rect 1390 3040 1405 3140
rect 1485 3040 1600 3140
rect 1390 3025 1600 3040
rect 1390 1640 1600 1655
rect 1390 1540 1405 1640
rect 1485 1540 1600 1640
rect 1390 1525 1600 1540
<< labels >>
rlabel metal3 625 1590 625 1590 7 bot
rlabel metal4 1600 1590 1600 1590 3 top
rlabel metal4 1600 3090 1600 3090 3 top
rlabel metal3 625 3090 625 3090 7 bot
<< end >>
