magic
tech sky130A
timestamp 1702791741
<< poly >>
rect -4525 8810 -4510 8820
rect -4980 8795 -4510 8810
rect -4815 8090 -4775 8100
rect -4815 8075 -4805 8090
rect -5010 8070 -4805 8075
rect -4785 8070 -4775 8090
rect -5010 8060 -4775 8070
<< polycont >>
rect -4805 8070 -4785 8090
<< locali >>
rect -4530 8735 -4090 8775
rect -4885 7385 -4865 8485
rect -4815 8090 -4775 8100
rect -4815 8070 -4805 8090
rect -4785 8080 -4775 8090
rect -4530 8080 -4510 8735
rect -4785 8070 -4510 8080
rect -4815 8060 -4510 8070
rect -5000 7365 -4865 7385
rect -5490 7080 -5450 7090
rect -5490 7030 -5480 7080
rect -5460 7030 -5450 7080
rect -5490 6935 -5450 7030
rect -5490 6925 -5410 6935
rect -5490 6905 -5480 6925
rect -5420 6905 -5410 6925
rect -5490 6895 -5410 6905
rect -5000 6620 -4980 7365
rect -5160 6600 -4980 6620
rect -4960 6865 -4915 6905
rect -4960 6345 -4940 6865
rect -5160 6325 -4940 6345
rect -5160 6050 -4905 6070
rect -5160 5775 -4945 5795
rect -5160 5500 -4985 5520
rect -5155 5225 -5025 5245
rect -5045 5150 -5025 5225
rect -5005 5195 -4985 5500
rect -4965 5240 -4945 5775
rect -4925 5705 -4905 6050
rect -4965 5220 -4915 5240
rect -5005 5175 -4955 5195
rect -5045 5130 -4995 5150
rect -5160 4950 -5035 4970
rect -5055 3540 -5035 4950
rect -5015 3585 -4995 5130
rect -4975 3630 -4955 5175
rect -4935 4105 -4915 5220
rect -4975 3610 -4890 3630
rect -5015 3565 -4945 3585
rect -5055 3520 -4990 3540
rect -6280 2185 -6250 3395
rect -6280 2150 -6185 2185
rect -6220 2060 -6185 2150
rect -6220 2050 -5935 2060
rect -6220 2030 -5995 2050
rect -5945 2030 -5935 2050
rect -6220 2020 -5935 2030
rect -5010 1990 -4990 3520
rect -4965 2035 -4945 3565
rect -4910 2540 -4890 3610
rect -4925 2500 -4890 2540
rect -4965 2015 -4865 2035
rect -5010 1970 -4945 1990
rect -6280 895 -6190 925
rect -6215 840 -6190 895
rect -6215 830 -6175 840
rect -6215 780 -6205 830
rect -6185 780 -6175 830
rect -6215 770 -6175 780
rect -4965 750 -4945 1970
rect -4885 1400 -4865 2015
rect -4925 1350 -4865 1400
rect -4965 720 -4810 750
rect 2745 680 2785 790
rect 2745 630 2755 680
rect 2775 630 2785 680
rect 2745 620 2785 630
<< viali >>
rect -5480 7030 -5460 7080
rect -5480 6905 -5420 6925
rect -5995 2030 -5945 2050
rect -6205 780 -6185 830
rect 2755 630 2775 680
<< metal1 >>
rect -4545 8735 -4395 8775
rect -4995 8690 -4530 8715
rect -4995 8115 -4870 8690
rect -4660 8675 -4530 8690
rect -4660 8670 -4595 8675
rect -6145 6845 -5685 7425
rect -4910 7250 -4870 8115
rect -5490 7205 -4870 7250
rect -5490 7080 -5450 7205
rect -5490 7030 -5480 7080
rect -5460 7030 -5450 7080
rect -5490 7020 -5450 7030
rect -5490 6925 -5410 6935
rect -5490 6905 -5480 6925
rect -5420 6905 -5410 6925
rect -5490 6880 -5410 6905
rect -5630 6830 -5160 6880
rect -6145 2305 -5685 2430
rect -6380 2275 -5685 2305
rect -6380 2090 -4810 2275
rect -5690 2085 -4810 2090
rect -6015 2050 -5865 2060
rect -6015 2030 -5995 2050
rect -5945 2030 -5865 2050
rect -6015 2020 -5865 2030
rect -6215 830 -6175 840
rect -6215 780 -6205 830
rect -6185 780 -6175 830
rect -6215 550 -6175 780
rect -5910 605 -5865 2020
rect 2810 785 2905 830
rect 2745 680 2785 690
rect 2745 630 2755 680
rect 2775 630 2785 680
rect 2745 605 2785 630
rect -5910 565 2785 605
rect 2860 550 2905 785
rect -6215 505 2905 550
use dac  dac_0 ~/VLSI_Sine_Gen/layout/dac
timestamp 1702787255
transform 1 0 -4510 0 1 7245
box -415 -6625 7355 1590
use filter  filter_0 ~/VLSI_Sine_Gen/layout/filter
timestamp 1702709769
transform -1 0 -5720 0 1 285
box 535 490 1685 3285
use register16  register16_0 ~/VLSI_Sine_Gen/layout/shift_register
timestamp 1702679440
transform 0 1 -6215 -1 0 6885
box -90 -15 4570 1140
use v_gen  v_gen_0 ~/VLSI_Sine_Gen/layout/v_gen
timestamp 1702787459
transform 1 0 -7075 0 1 7375
box -35 -10 2120 1435
<< end >>
