magic
tech sky130A
timestamp 1702790376
<< psubdiff >>
rect 715 2940 865 2955
rect 715 2910 730 2940
rect 850 2910 865 2940
rect 715 2895 865 2910
rect 810 2800 870 2815
rect 810 2680 825 2800
rect 855 2680 870 2800
rect 810 2665 870 2680
rect 620 1920 680 1935
rect 620 1800 635 1920
rect 665 1800 680 1920
rect 620 1785 680 1800
rect 630 1110 690 1125
rect 630 990 645 1110
rect 675 990 690 1110
rect 630 975 690 990
rect 1665 800 1815 815
rect 1665 770 1680 800
rect 1800 770 1815 800
rect 1665 755 1815 770
<< psubdiffcont >>
rect 730 2910 850 2940
rect 825 2680 855 2800
rect 635 1800 665 1920
rect 645 990 675 1110
rect 1680 770 1800 800
<< xpolycontact >>
rect 930 2945 1150 2980
rect 1500 2945 1720 2980
rect 930 2885 1150 2920
rect 1500 2885 1720 2920
rect 930 2770 1150 2805
rect 1500 2770 1720 2805
rect 930 2665 1150 2700
rect 1500 2665 1720 2700
rect 600 1700 820 1735
rect 1170 1700 1390 1735
rect 545 1325 580 1545
rect 545 755 580 975
rect 780 810 1000 845
rect 1350 810 1570 845
rect 780 750 1000 785
rect 1350 750 1570 785
<< xpolyres >>
rect 1150 2945 1500 2980
rect 1150 2885 1500 2920
rect 1150 2770 1500 2805
rect 1150 2665 1500 2700
rect 820 1700 1170 1735
rect 545 975 580 1325
rect 1000 810 1350 845
rect 1000 750 1350 785
<< locali >>
rect 720 2940 860 2950
rect 720 2910 730 2940
rect 850 2910 860 2940
rect 720 2900 860 2910
rect 1720 2965 1800 2980
rect 1720 2945 1755 2965
rect 930 2920 1150 2945
rect 1500 2865 1720 2885
rect 535 2840 1720 2865
rect 1740 2860 1755 2945
rect 1785 2860 1800 2965
rect 1740 2845 1800 2860
rect 815 2800 865 2810
rect 1500 2805 1720 2840
rect 815 2680 825 2800
rect 855 2680 865 2800
rect 815 2670 865 2680
rect 930 2755 1150 2770
rect 930 2745 1080 2755
rect 930 2715 945 2745
rect 1065 2715 1080 2745
rect 930 2700 1080 2715
rect 1720 2665 1835 2700
rect 1795 2655 1835 2665
rect 1795 2595 1875 2655
rect 1795 2495 1810 2595
rect 1860 2495 1875 2595
rect 1795 2480 1875 2495
rect 1795 2000 1875 2015
rect 625 1920 675 1930
rect 625 1800 635 1920
rect 665 1800 675 1920
rect 625 1790 675 1800
rect 1795 1900 1810 2000
rect 1860 1900 1875 2000
rect 1795 1735 1875 1900
rect 545 1700 600 1735
rect 1390 1700 1885 1735
rect 545 1680 580 1700
rect 545 1665 625 1680
rect 545 1565 560 1665
rect 610 1565 625 1665
rect 545 1550 625 1565
rect 1800 1640 1880 1655
rect 545 1545 580 1550
rect 1800 1540 1815 1640
rect 1865 1540 1880 1640
rect 1800 1525 1880 1540
rect 635 1110 685 1120
rect 635 990 645 1110
rect 675 990 685 1110
rect 635 980 685 990
rect 535 755 545 845
rect 580 810 780 845
rect 580 755 595 810
rect 650 785 1000 790
rect 650 780 780 785
rect 650 750 665 780
rect 765 750 780 780
rect 1350 785 1570 810
rect 1670 800 1810 810
rect 1670 770 1680 800
rect 1800 770 1810 800
rect 1670 760 1810 770
rect 650 740 1000 750
<< viali >>
rect 730 2910 850 2940
rect 1755 2860 1785 2965
rect 825 2680 855 2800
rect 945 2715 1065 2745
rect 1810 2495 1860 2595
rect 635 1800 665 1920
rect 1810 1900 1860 2000
rect 560 1565 610 1665
rect 1815 1540 1865 1640
rect 645 990 675 1110
rect 665 750 765 780
rect 1680 770 1800 800
<< metal1 >>
rect 650 2940 910 2980
rect 650 2910 730 2940
rect 850 2910 910 2940
rect 650 2875 910 2910
rect 1740 2965 1845 2980
rect 1740 2875 1755 2965
rect 650 2860 1755 2875
rect 1785 2860 1845 2965
rect 650 2825 1845 2860
rect 650 2800 910 2825
rect 650 2680 825 2800
rect 855 2680 910 2800
rect 930 2745 1080 2760
rect 930 2715 945 2745
rect 1065 2715 1080 2745
rect 930 2700 1080 2715
rect 650 2645 910 2680
rect 650 1975 690 2645
rect 1795 2595 1875 2610
rect 1795 2495 1810 2595
rect 1860 2495 1875 2595
rect 1795 2480 1875 2495
rect 600 1920 690 1975
rect 600 1800 635 1920
rect 665 1800 690 1920
rect 1795 2000 1875 2015
rect 1795 1900 1810 2000
rect 1860 1900 1875 2000
rect 1795 1885 1875 1900
rect 600 1770 690 1800
rect 545 1665 625 1680
rect 545 1565 560 1665
rect 610 1565 625 1665
rect 545 1550 625 1565
rect 650 1520 690 1770
rect 1800 1640 1880 1655
rect 1800 1540 1815 1640
rect 1865 1540 1880 1640
rect 1800 1525 1880 1540
rect 630 1110 690 1520
rect 630 990 645 1110
rect 675 990 690 1110
rect 630 800 690 990
rect 1625 800 1885 850
rect 630 780 1680 800
rect 630 750 665 780
rect 765 770 1680 780
rect 1800 770 1885 800
rect 765 750 1885 770
rect 630 740 1885 750
<< via1 >>
rect 945 2715 1065 2745
rect 1810 2495 1860 2595
rect 1810 1900 1860 2000
rect 560 1565 610 1665
rect 1815 1540 1865 1640
<< metal2 >>
rect 930 2745 1080 2760
rect 930 2715 945 2745
rect 1065 2730 1080 2745
rect 1065 2715 1775 2730
rect 930 2700 1775 2715
rect 545 1665 625 1680
rect 545 1565 560 1665
rect 610 1565 625 1665
rect 545 1550 625 1565
rect 1745 1655 1775 2700
rect 1795 2595 1875 2610
rect 1795 2495 1810 2595
rect 1860 2495 1875 2595
rect 1795 2480 1875 2495
rect 1795 2000 1875 2015
rect 1795 1900 1810 2000
rect 1860 1900 1875 2000
rect 1795 1885 1875 1900
rect 1745 1640 1880 1655
rect 1745 1540 1815 1640
rect 1865 1540 1880 1640
rect 1745 1525 1880 1540
<< via2 >>
rect 560 1565 610 1665
rect 1810 2495 1860 2595
rect 1810 1900 1860 2000
rect 1815 1540 1865 1640
<< metal3 >>
rect 690 2015 1730 2645
rect 1795 2595 1875 2610
rect 1795 2495 1810 2595
rect 1860 2495 1875 2595
rect 1795 2480 1875 2495
rect 690 2000 1875 2015
rect 690 1900 1810 2000
rect 1860 1900 1875 2000
rect 690 1885 1875 1900
rect 690 1805 1730 1885
rect 700 1680 1730 1685
rect 545 1665 1730 1680
rect 545 1565 560 1665
rect 610 1565 1730 1665
rect 545 1550 1730 1565
rect 700 855 1730 1550
rect 1800 1640 1880 1655
rect 1800 1540 1815 1640
rect 1865 1540 1880 1640
rect 1800 1525 1880 1540
<< via3 >>
rect 1810 2495 1860 2595
rect 1815 1540 1865 1640
<< mimcap >>
rect 710 2595 1710 2625
rect 710 2495 1600 2595
rect 1680 2495 1710 2595
rect 710 1825 1710 2495
rect 715 1640 1715 1670
rect 715 1540 1605 1640
rect 1685 1540 1715 1640
rect 715 870 1715 1540
<< mimcapcontact >>
rect 1600 2495 1680 2595
rect 1605 1540 1685 1640
<< metal4 >>
rect 1585 2595 1875 2610
rect 1585 2495 1600 2595
rect 1680 2495 1810 2595
rect 1860 2495 1875 2595
rect 1585 2480 1875 2495
rect 1590 1640 1880 1655
rect 1590 1540 1605 1640
rect 1685 1540 1815 1640
rect 1865 1540 1880 1640
rect 1590 1525 1880 1540
<< labels >>
rlabel locali 1885 1720 1885 1720 3 Vout-
rlabel locali 535 825 535 825 7 Viout-
rlabel locali 535 2855 535 2855 7 Viout+
rlabel xpolycontact 1685 2685 1685 2685 3 Vout+
rlabel metal1 1885 790 1885 790 3 VN
<< end >>
