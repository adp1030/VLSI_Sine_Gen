magic
tech sky130A
timestamp 1702715363
<< poly >>
rect 8975 6870 9115 6880
rect 8975 6850 8985 6870
rect 9005 6860 9085 6870
rect 9005 6850 9015 6860
rect 8975 6840 9015 6850
rect 9075 6850 9085 6860
rect 9105 6850 9115 6870
rect 9075 6840 9115 6850
rect 9855 5895 10155 5915
rect 9855 5855 9875 5895
rect 9915 5855 10095 5895
rect 10135 5855 10155 5895
rect 9855 5835 10155 5855
<< polycont >>
rect 8985 6850 9005 6870
rect 9085 6850 9105 6870
rect 9875 5855 9915 5895
rect 10095 5855 10135 5895
<< locali >>
rect 9035 6900 9925 6920
rect 8975 6870 9015 6880
rect 8975 6850 8985 6870
rect 9005 6850 9015 6870
rect 8975 6840 9015 6850
rect 8995 6825 9015 6835
rect 9035 6790 9055 6900
rect 9075 6870 9920 6880
rect 9075 6850 9085 6870
rect 9105 6860 9920 6870
rect 9105 6850 9115 6860
rect 9075 6840 9115 6850
rect 9805 6775 9895 6795
rect 9310 4210 9415 4220
rect 9310 4190 9320 4210
rect 9405 4190 9415 4210
rect 9310 4095 9415 4190
rect 9805 4140 9825 6775
rect 9855 5895 9935 5915
rect 9855 5855 9875 5895
rect 9915 5855 9935 5895
rect 9855 5835 9935 5855
rect 10075 5895 10155 5915
rect 10075 5855 10095 5895
rect 10135 5855 10155 5895
rect 10075 5835 10155 5855
rect 9310 4075 9320 4095
rect 9405 4075 9415 4095
rect 9310 4065 9415 4075
rect 9785 4120 9825 4140
rect 9845 5665 9890 5685
rect 9785 3805 9805 4120
rect 9845 4100 9865 5665
rect 9635 3785 9805 3805
rect 9825 4080 9865 4100
rect 9825 3530 9845 4080
rect 9595 3510 9845 3530
rect 9865 3740 9910 3760
rect 9865 3255 9885 3740
rect 9635 3235 9885 3255
rect 9570 2960 9855 2980
rect 9570 2685 9815 2705
rect 9600 2410 9775 2430
rect 9550 2135 9735 2155
rect 9715 -2970 9735 2135
rect 9755 -2015 9775 2410
rect 9795 -90 9815 2685
rect 9835 1835 9855 2960
rect 18915 2030 18955 2040
rect 18915 1980 18925 2030
rect 18945 1980 18955 2030
rect 9835 1815 9900 1835
rect 18915 1810 18955 1980
rect 20340 2030 20380 2040
rect 20340 1980 20350 2030
rect 20370 1980 20380 2030
rect 20340 1970 20380 1980
rect 18915 1785 19005 1810
rect 9970 900 9975 920
rect 9795 -110 9900 -90
rect 18875 -665 19000 -655
rect 18875 -715 18885 -665
rect 18905 -690 19000 -665
rect 18905 -715 18915 -690
rect 18875 -725 18915 -715
rect 20300 -850 20340 -840
rect 20300 -900 20310 -850
rect 20330 -900 20340 -850
rect 20300 -910 20340 -900
rect 9755 -2035 9895 -2015
rect 20320 -2950 20340 -910
rect 20300 -2970 20340 -2950
rect 9715 -2990 9895 -2970
rect 20360 -2990 20380 1970
rect 20280 -3010 20380 -2990
<< viali >>
rect 9320 4190 9405 4210
rect 9875 5855 9915 5895
rect 10095 5855 10135 5895
rect 9320 4075 9405 4095
rect 18925 1980 18945 2030
rect 20350 1980 20370 2030
rect 18885 -715 18905 -665
rect 20310 -900 20330 -850
<< metal1 >>
rect 9690 5895 9940 5915
rect 9690 5855 9875 5895
rect 9915 5855 9940 5895
rect 9690 5835 9940 5855
rect 10075 5895 10350 5915
rect 10075 5855 10095 5895
rect 10135 5855 10350 5895
rect 10075 5835 10350 5855
rect 8370 4580 8970 4600
rect 9090 4580 9690 4595
rect 8665 4065 8750 4580
rect 9310 4210 9415 4580
rect 10280 4450 10350 5015
rect 9310 4190 9320 4210
rect 9405 4190 9415 4210
rect 9310 4180 9415 4190
rect 9310 4095 9415 4105
rect 9310 4075 9320 4095
rect 9405 4075 9415 4095
rect 9310 4065 9415 4075
rect 8665 4045 9125 4065
rect 9180 4030 9650 4065
rect 10275 2530 10345 3095
rect 18915 2030 20380 2040
rect 18915 1980 18925 2030
rect 18945 2010 20350 2030
rect 18945 1980 18955 2010
rect 18915 1970 18955 1980
rect 20340 1980 20350 2010
rect 20370 1980 20380 2030
rect 20340 1970 20380 1980
rect 10275 590 10345 1155
rect 8665 -405 9125 -375
rect 8900 -2840 8945 -405
rect 18875 -665 18915 -655
rect 18875 -715 18885 -665
rect 18905 -715 18915 -665
rect 10275 -1335 10345 -770
rect 18875 -840 18915 -715
rect 19925 -810 20390 -735
rect 18875 -850 20340 -840
rect 18875 -875 20310 -850
rect 20300 -900 20310 -875
rect 20330 -900 20340 -850
rect 20300 -910 20340 -900
rect 8900 -2845 9250 -2840
rect 20360 -2845 20390 -810
rect 8900 -2885 20390 -2845
rect 8905 -2890 20390 -2885
use dac_v2  dac_v2_0 ~/VLSI_Sine_Gen/layout/dac
timestamp 1702516191
transform 1 0 10275 0 1 6855
box -400 -9865 10045 65
use filter  filter_0 ~/VLSI_Sine_Gen/layout/filter
timestamp 1702709769
transform 1 0 18405 0 1 -1300
box 535 490 1685 3285
use register16  register16_0 ~/VLSI_Sine_Gen/layout/shift_register
timestamp 1702679440
transform 0 1 8595 -1 0 4070
box -90 -15 4570 1140
use v_gen  v_gen_0 ~/VLSI_Sine_Gen/layout/bias_gen
timestamp 1702521636
transform 0 1 8340 1 0 4700
box -120 -55 2140 1445
<< end >>
