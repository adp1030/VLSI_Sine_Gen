* NGSPICE file created from dac_v2.ext - technology: sky130A

.subckt dac_unit Vphi Vphi_b Vbp Vcp Viun Viup VP
X0 a_1440_150# Vcp a_1070_1810# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X1 VP Vbp a_100_150# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X2 a_1440_150# Vbp VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X3 a_300_150# Vcp a_100_150# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X4 Viup Vphi_b a_300_150# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=3 ps=13 w=6 l=0.5
X5 a_1070_1810# Vphi_b Viup VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=3 ps=13 w=6 l=0.5
X6 VP VP a_1440_150# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X7 a_100_150# VP VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X8 a_1070_1810# Vphi Viun VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X9 a_100_150# VP VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X10 Viun Vphi a_300_150# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X11 VP VP a_1440_150# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
.ends

.subckt inverter A Y VP VN
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
.ends

Xdac_unit_4 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_5 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_6 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xinverter_0 Vphi7 inverter_0/Y inverter_7/VP VSUBS inverter
Xinverter_1 Vphi2 inverter_1/Y inverter_7/VP VSUBS inverter
Xdac_unit_7 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_8 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xinverter_2 Vphi3 inverter_2/Y inverter_7/VP VSUBS inverter
Xinverter_3 Vphi4 inverter_3/Y inverter_7/VP VSUBS inverter
Xdac_unit_9 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xinverter_4 Vphi5 inverter_4/Y inverter_7/VP VSUBS inverter
Xinverter_5 Vphi6 inverter_5/Y inverter_7/VP VSUBS inverter
Xinverter_7 Vphi1 inverter_7/Y inverter_7/VP VSUBS inverter
Xdac_unit_40 Vphi1 inverter_7/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_41 Vphi1 inverter_7/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_30 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_42 Vphi1 inverter_7/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_20 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_31 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_10 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_21 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_32 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_11 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_22 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_33 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_12 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_23 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_34 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_14 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_13 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_25 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_24 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_36 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_35 Vphi6 inverter_5/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_15 Vphi3 inverter_2/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_26 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_16 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_27 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_17 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_28 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_18 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_29 Vphi5 inverter_4/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_19 Vphi4 inverter_3/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_0 Vphi7 inverter_0/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_1 Vphi7 inverter_0/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_2 Vphi7 inverter_0/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit
Xdac_unit_3 Vphi2 inverter_1/Y Vbp Vcp Viout- Viout+ inverter_7/VP dac_unit

