** sch_path: /home/madvlsi/VLSI_Sine_Gen/simulation/filter/cap.sch
**.subckt cap
XC3 top bot sky130_fd_pr__cap_mim_m3_1 W=10 L=8 MF=1 m=1
XC1 top bot sky130_fd_pr__cap_mim_m3_1 W=10 L=8 MF=1 m=1
**.ends
.end
