magic
tech sky130A
timestamp 1702620399
<< nwell >>
rect 4835 105 4950 1460
rect 5635 -1495 5755 -140
rect 5635 -4700 5765 -3345
rect 4835 -6305 4975 -4950
<< poly >>
rect 5330 -20 5370 -10
rect 5330 -40 5340 -20
rect 5360 -25 5370 -20
rect 6130 -20 6170 -10
rect 6130 -25 6140 -20
rect 5360 -40 6140 -25
rect 6160 -40 6170 -20
rect 5330 -50 6170 -40
rect 5330 -6430 5370 -6420
rect 5330 -6450 5340 -6430
rect 5360 -6435 5370 -6430
rect 6130 -6430 6170 -6420
rect 6130 -6435 6140 -6430
rect 5360 -6450 6140 -6435
rect 6160 -6450 6170 -6430
rect 5330 -6460 6170 -6450
<< polycont >>
rect 5340 -40 5360 -20
rect 6140 -40 6160 -20
rect 5340 -6450 5360 -6430
rect 6140 -6450 6160 -6430
<< locali >>
rect -70 90 0 100
rect -70 70 -60 90
rect -10 70 0 90
rect -70 60 0 70
rect 225 -65 260 45
rect 430 -10 460 45
rect 430 -20 500 -10
rect 430 -40 440 -20
rect 490 -40 500 -20
rect 430 -50 500 -40
rect 1025 -65 1060 45
rect 1230 -10 1260 45
rect 1230 -20 1300 -10
rect 1230 -40 1240 -20
rect 1290 -40 1300 -20
rect 1230 -50 1300 -40
rect 1825 -65 1860 45
rect 2030 -10 2060 45
rect 2030 -20 2100 -10
rect 2030 -40 2040 -20
rect 2090 -40 2100 -20
rect 2030 -50 2100 -40
rect 2625 -65 2660 45
rect 2830 -10 2860 45
rect 2830 -20 2900 -10
rect 2830 -40 2840 -20
rect 2890 -40 2900 -20
rect 2830 -50 2900 -40
rect 3425 -65 3460 45
rect 3630 -10 3660 45
rect 3630 -20 3700 -10
rect 3630 -40 3640 -20
rect 3690 -40 3700 -20
rect 3630 -50 3700 -40
rect 4225 -65 4260 45
rect 4430 -10 4460 45
rect 4430 -20 4500 -10
rect 4430 -40 4440 -20
rect 4490 -40 4500 -20
rect 4430 -50 4500 -40
rect 225 -75 295 -65
rect 225 -95 235 -75
rect 285 -95 295 -75
rect 225 -105 295 -95
rect 1025 -75 1095 -65
rect 1025 -95 1035 -75
rect 1085 -95 1095 -75
rect 1025 -105 1095 -95
rect 1825 -75 1895 -65
rect 1825 -95 1835 -75
rect 1885 -95 1895 -75
rect 1825 -105 1895 -95
rect 2625 -75 2695 -65
rect 2625 -95 2635 -75
rect 2685 -95 2695 -75
rect 2625 -105 2695 -95
rect 3425 -75 3495 -65
rect 3425 -95 3435 -75
rect 3485 -95 3495 -75
rect 3425 -105 3495 -95
rect 4225 -75 4295 -65
rect 4225 -95 4235 -75
rect 4285 -95 4295 -75
rect 4225 -105 4295 -95
rect 5130 -80 5165 15
rect 5335 -10 5365 5
rect 5330 -20 5370 -10
rect 5330 -40 5340 -20
rect 5360 -40 5370 -20
rect 5330 -50 5370 -40
rect 5930 -80 5965 15
rect 6135 -10 6165 50
rect 6130 -20 6170 -10
rect 6130 -40 6140 -20
rect 6160 -25 6170 -20
rect 6160 -40 6595 -25
rect 6130 -50 6595 -40
rect 5130 -105 6595 -80
rect -70 -1510 0 -1500
rect -70 -1530 -60 -1510
rect -10 -1530 0 -1510
rect -70 -1540 0 -1530
rect 225 -1665 260 -1555
rect 430 -1610 460 -1555
rect 430 -1620 500 -1610
rect 430 -1640 440 -1620
rect 490 -1640 500 -1620
rect 430 -1650 500 -1640
rect 1025 -1665 1060 -1555
rect 1230 -1610 1260 -1555
rect 1230 -1620 1300 -1610
rect 1230 -1640 1240 -1620
rect 1290 -1640 1300 -1620
rect 1230 -1650 1300 -1640
rect 1825 -1665 1860 -1555
rect 2030 -1610 2060 -1555
rect 2030 -1620 2100 -1610
rect 2030 -1640 2040 -1620
rect 2090 -1640 2100 -1620
rect 2030 -1650 2100 -1640
rect 2625 -1665 2660 -1555
rect 2830 -1610 2860 -1555
rect 2830 -1620 2900 -1610
rect 2830 -1640 2840 -1620
rect 2890 -1640 2900 -1620
rect 2830 -1650 2900 -1640
rect 3425 -1665 3460 -1555
rect 3630 -1610 3660 -1555
rect 3630 -1620 3700 -1610
rect 3630 -1640 3640 -1620
rect 3690 -1640 3700 -1620
rect 3630 -1650 3700 -1640
rect 4225 -1665 4260 -1555
rect 4430 -1610 4460 -1555
rect 4430 -1620 4500 -1610
rect 4430 -1640 4440 -1620
rect 4490 -1640 4500 -1620
rect 4430 -1650 4500 -1640
rect 5025 -1665 5060 -1555
rect 5230 -1610 5260 -1555
rect 5230 -1620 5300 -1610
rect 5230 -1640 5240 -1620
rect 5290 -1640 5300 -1620
rect 5230 -1650 5300 -1640
rect 225 -1675 295 -1665
rect 225 -1695 235 -1675
rect 285 -1695 295 -1675
rect 225 -1705 295 -1695
rect 1025 -1675 1095 -1665
rect 1025 -1695 1035 -1675
rect 1085 -1695 1095 -1675
rect 1025 -1705 1095 -1695
rect 1825 -1675 1895 -1665
rect 1825 -1695 1835 -1675
rect 1885 -1695 1895 -1675
rect 1825 -1705 1895 -1695
rect 2625 -1675 2695 -1665
rect 2625 -1695 2635 -1675
rect 2685 -1695 2695 -1675
rect 2625 -1705 2695 -1695
rect 3425 -1675 3495 -1665
rect 3425 -1695 3435 -1675
rect 3485 -1695 3495 -1675
rect 3425 -1705 3495 -1695
rect 4225 -1675 4295 -1665
rect 4225 -1695 4235 -1675
rect 4285 -1695 4295 -1675
rect 4225 -1705 4295 -1695
rect 5025 -1675 5095 -1665
rect 5025 -1695 5035 -1675
rect 5085 -1695 5095 -1675
rect 5025 -1705 5095 -1695
rect -70 -3110 0 -3100
rect -70 -3130 -60 -3110
rect -10 -3130 0 -3110
rect -70 -3140 0 -3130
rect 225 -3265 260 -3155
rect 430 -3210 460 -3155
rect 430 -3220 500 -3210
rect 430 -3240 440 -3220
rect 490 -3240 500 -3220
rect 430 -3250 500 -3240
rect 1025 -3265 1060 -3155
rect 1230 -3210 1260 -3155
rect 1230 -3220 1300 -3210
rect 1230 -3240 1240 -3220
rect 1290 -3240 1300 -3220
rect 1230 -3250 1300 -3240
rect 1825 -3265 1860 -3155
rect 2030 -3210 2060 -3155
rect 2030 -3220 2100 -3210
rect 2030 -3240 2040 -3220
rect 2090 -3240 2100 -3220
rect 2030 -3250 2100 -3240
rect 2625 -3265 2660 -3155
rect 2830 -3210 2860 -3155
rect 2830 -3220 2900 -3210
rect 2830 -3240 2840 -3220
rect 2890 -3240 2900 -3220
rect 2830 -3250 2900 -3240
rect 3425 -3265 3460 -3155
rect 3630 -3210 3660 -3155
rect 3630 -3220 3700 -3210
rect 3630 -3240 3640 -3220
rect 3690 -3240 3700 -3220
rect 3630 -3250 3700 -3240
rect 4225 -3265 4260 -3155
rect 4430 -3210 4460 -3155
rect 4430 -3220 4500 -3210
rect 4430 -3240 4440 -3220
rect 4490 -3240 4500 -3220
rect 4430 -3250 4500 -3240
rect 5025 -3265 5060 -3155
rect 5230 -3210 5260 -3155
rect 5230 -3220 5300 -3210
rect 5230 -3240 5240 -3220
rect 5290 -3240 5300 -3220
rect 5230 -3250 5300 -3240
rect 5825 -3265 5860 -3155
rect 6030 -3210 6060 -3155
rect 6030 -3220 6100 -3210
rect 6030 -3240 6040 -3220
rect 6090 -3240 6100 -3220
rect 6030 -3250 6100 -3240
rect 225 -3275 295 -3265
rect 225 -3295 235 -3275
rect 285 -3295 295 -3275
rect 225 -3305 295 -3295
rect 1025 -3275 1095 -3265
rect 1025 -3295 1035 -3275
rect 1085 -3295 1095 -3275
rect 1025 -3305 1095 -3295
rect 1825 -3275 1895 -3265
rect 1825 -3295 1835 -3275
rect 1885 -3295 1895 -3275
rect 1825 -3305 1895 -3295
rect 2625 -3275 2695 -3265
rect 2625 -3295 2635 -3275
rect 2685 -3295 2695 -3275
rect 2625 -3305 2695 -3295
rect 3425 -3275 3495 -3265
rect 3425 -3295 3435 -3275
rect 3485 -3295 3495 -3275
rect 3425 -3305 3495 -3295
rect 4225 -3275 4295 -3265
rect 4225 -3295 4235 -3275
rect 4285 -3295 4295 -3275
rect 4225 -3305 4295 -3295
rect 5025 -3275 5095 -3265
rect 5025 -3295 5035 -3275
rect 5085 -3295 5095 -3275
rect 5025 -3305 5095 -3295
rect 5825 -3275 5895 -3265
rect 5825 -3295 5835 -3275
rect 5885 -3295 5895 -3275
rect 5825 -3305 5895 -3295
rect -70 -4715 0 -4705
rect -70 -4735 -60 -4715
rect -10 -4735 0 -4715
rect -70 -4745 0 -4735
rect 225 -4870 260 -4760
rect 430 -4815 460 -4760
rect 430 -4825 500 -4815
rect 430 -4845 440 -4825
rect 490 -4845 500 -4825
rect 430 -4855 500 -4845
rect 1025 -4870 1060 -4760
rect 1230 -4815 1260 -4760
rect 1230 -4825 1300 -4815
rect 1230 -4845 1240 -4825
rect 1290 -4845 1300 -4825
rect 1230 -4855 1300 -4845
rect 1825 -4870 1860 -4760
rect 2030 -4815 2060 -4760
rect 2030 -4825 2100 -4815
rect 2030 -4845 2040 -4825
rect 2090 -4845 2100 -4825
rect 2030 -4855 2100 -4845
rect 2625 -4870 2660 -4760
rect 2830 -4815 2860 -4760
rect 2830 -4825 2900 -4815
rect 2830 -4845 2840 -4825
rect 2890 -4845 2900 -4825
rect 2830 -4855 2900 -4845
rect 3425 -4870 3460 -4760
rect 3630 -4815 3660 -4760
rect 3630 -4825 3700 -4815
rect 3630 -4845 3640 -4825
rect 3690 -4845 3700 -4825
rect 3630 -4855 3700 -4845
rect 4225 -4870 4260 -4760
rect 4430 -4815 4460 -4760
rect 4430 -4825 4500 -4815
rect 4430 -4845 4440 -4825
rect 4490 -4845 4500 -4825
rect 4430 -4855 4500 -4845
rect 5025 -4870 5060 -4760
rect 5230 -4815 5260 -4760
rect 5230 -4825 5300 -4815
rect 5230 -4845 5240 -4825
rect 5290 -4845 5300 -4825
rect 5230 -4855 5300 -4845
rect 225 -4880 295 -4870
rect 225 -4900 235 -4880
rect 285 -4900 295 -4880
rect 225 -4910 295 -4900
rect 1025 -4880 1095 -4870
rect 1025 -4900 1035 -4880
rect 1085 -4900 1095 -4880
rect 1025 -4910 1095 -4900
rect 1825 -4880 1895 -4870
rect 1825 -4900 1835 -4880
rect 1885 -4900 1895 -4880
rect 1825 -4910 1895 -4900
rect 2625 -4880 2695 -4870
rect 2625 -4900 2635 -4880
rect 2685 -4900 2695 -4880
rect 2625 -4910 2695 -4900
rect 3425 -4880 3495 -4870
rect 3425 -4900 3435 -4880
rect 3485 -4900 3495 -4880
rect 3425 -4910 3495 -4900
rect 4225 -4880 4295 -4870
rect 4225 -4900 4235 -4880
rect 4285 -4900 4295 -4880
rect 4225 -4910 4295 -4900
rect 5025 -4880 5095 -4870
rect 5025 -4900 5035 -4880
rect 5085 -4900 5095 -4880
rect 5025 -4910 5095 -4900
rect -70 -6320 0 -6310
rect -70 -6340 -60 -6320
rect -10 -6340 0 -6320
rect -70 -6350 0 -6340
rect 225 -6475 260 -6365
rect 430 -6420 460 -6365
rect 430 -6430 500 -6420
rect 430 -6450 440 -6430
rect 490 -6450 500 -6430
rect 430 -6460 500 -6450
rect 1025 -6475 1060 -6365
rect 1230 -6420 1260 -6365
rect 1230 -6430 1300 -6420
rect 1230 -6450 1240 -6430
rect 1290 -6450 1300 -6430
rect 1230 -6460 1300 -6450
rect 1825 -6475 1860 -6365
rect 2030 -6420 2060 -6365
rect 2030 -6430 2100 -6420
rect 2030 -6450 2040 -6430
rect 2090 -6450 2100 -6430
rect 2030 -6460 2100 -6450
rect 2625 -6475 2660 -6365
rect 2830 -6420 2860 -6365
rect 2830 -6430 2900 -6420
rect 2830 -6450 2840 -6430
rect 2890 -6450 2900 -6430
rect 2830 -6460 2900 -6450
rect 3425 -6475 3460 -6365
rect 3630 -6420 3660 -6365
rect 3630 -6430 3700 -6420
rect 3630 -6450 3640 -6430
rect 3690 -6450 3700 -6430
rect 3630 -6460 3700 -6450
rect 4225 -6475 4260 -6365
rect 4430 -6420 4460 -6365
rect 4430 -6430 4500 -6420
rect 4430 -6450 4440 -6430
rect 4490 -6450 4500 -6430
rect 4430 -6460 4500 -6450
rect 225 -6485 295 -6475
rect 225 -6505 235 -6485
rect 285 -6505 295 -6485
rect 225 -6515 295 -6505
rect 1025 -6485 1095 -6475
rect 1025 -6505 1035 -6485
rect 1085 -6505 1095 -6485
rect 1025 -6515 1095 -6505
rect 1825 -6485 1895 -6475
rect 1825 -6505 1835 -6485
rect 1885 -6505 1895 -6485
rect 1825 -6515 1895 -6505
rect 2625 -6485 2695 -6475
rect 2625 -6505 2635 -6485
rect 2685 -6505 2695 -6485
rect 2625 -6515 2695 -6505
rect 3425 -6485 3495 -6475
rect 3425 -6505 3435 -6485
rect 3485 -6505 3495 -6485
rect 3425 -6515 3495 -6505
rect 4225 -6485 4295 -6475
rect 4225 -6505 4235 -6485
rect 4285 -6505 4295 -6485
rect 4225 -6515 4295 -6505
rect 5130 -6490 5165 -6395
rect 5335 -6420 5365 -6405
rect 5330 -6430 5370 -6420
rect 5330 -6450 5340 -6430
rect 5360 -6450 5370 -6430
rect 5330 -6460 5370 -6450
rect 5930 -6490 5965 -6395
rect 6135 -6420 6165 -6360
rect 6130 -6430 6170 -6420
rect 6130 -6450 6140 -6430
rect 6160 -6435 6170 -6430
rect 6160 -6450 6595 -6435
rect 6130 -6460 6595 -6450
rect 5130 -6515 6595 -6490
<< viali >>
rect -60 70 -10 90
rect 440 -40 490 -20
rect 1240 -40 1290 -20
rect 2040 -40 2090 -20
rect 2840 -40 2890 -20
rect 3640 -40 3690 -20
rect 4440 -40 4490 -20
rect 235 -95 285 -75
rect 1035 -95 1085 -75
rect 1835 -95 1885 -75
rect 2635 -95 2685 -75
rect 3435 -95 3485 -75
rect 4235 -95 4285 -75
rect -60 -1530 -10 -1510
rect 440 -1640 490 -1620
rect 1240 -1640 1290 -1620
rect 2040 -1640 2090 -1620
rect 2840 -1640 2890 -1620
rect 3640 -1640 3690 -1620
rect 4440 -1640 4490 -1620
rect 5240 -1640 5290 -1620
rect 235 -1695 285 -1675
rect 1035 -1695 1085 -1675
rect 1835 -1695 1885 -1675
rect 2635 -1695 2685 -1675
rect 3435 -1695 3485 -1675
rect 4235 -1695 4285 -1675
rect 5035 -1695 5085 -1675
rect -60 -3130 -10 -3110
rect 440 -3240 490 -3220
rect 1240 -3240 1290 -3220
rect 2040 -3240 2090 -3220
rect 2840 -3240 2890 -3220
rect 3640 -3240 3690 -3220
rect 4440 -3240 4490 -3220
rect 5240 -3240 5290 -3220
rect 6040 -3240 6090 -3220
rect 235 -3295 285 -3275
rect 1035 -3295 1085 -3275
rect 1835 -3295 1885 -3275
rect 2635 -3295 2685 -3275
rect 3435 -3295 3485 -3275
rect 4235 -3295 4285 -3275
rect 5035 -3295 5085 -3275
rect 5835 -3295 5885 -3275
rect -60 -4735 -10 -4715
rect 440 -4845 490 -4825
rect 1240 -4845 1290 -4825
rect 2040 -4845 2090 -4825
rect 2840 -4845 2890 -4825
rect 3640 -4845 3690 -4825
rect 4440 -4845 4490 -4825
rect 5240 -4845 5290 -4825
rect 235 -4900 285 -4880
rect 1035 -4900 1085 -4880
rect 1835 -4900 1885 -4880
rect 2635 -4900 2685 -4880
rect 3435 -4900 3485 -4880
rect 4235 -4900 4285 -4880
rect 5035 -4900 5085 -4880
rect -60 -6340 -10 -6320
rect 440 -6450 490 -6430
rect 1240 -6450 1290 -6430
rect 2040 -6450 2090 -6430
rect 2840 -6450 2890 -6430
rect 3640 -6450 3690 -6430
rect 4440 -6450 4490 -6430
rect 235 -6505 285 -6485
rect 1035 -6505 1085 -6485
rect 1835 -6505 1885 -6485
rect 2635 -6505 2685 -6485
rect 3435 -6505 3485 -6485
rect 4235 -6505 4285 -6485
<< metal1 >>
rect 4845 135 4945 1430
rect -70 90 70 100
rect -70 70 -60 90
rect -10 70 70 90
rect -70 60 70 70
rect 6595 60 6620 100
rect -70 5 70 45
rect 6595 5 6620 45
rect 430 -20 6595 -10
rect 430 -40 440 -20
rect 490 -40 1240 -20
rect 1290 -40 2040 -20
rect 2090 -40 2840 -20
rect 2890 -40 3640 -20
rect 3690 -40 4440 -20
rect 4490 -40 6595 -20
rect 430 -50 6595 -40
rect 225 -75 6595 -65
rect 225 -95 235 -75
rect 285 -95 1035 -75
rect 1085 -95 1835 -75
rect 1885 -95 2635 -75
rect 2685 -95 3435 -75
rect 3485 -95 4235 -75
rect 4285 -95 6595 -75
rect 225 -105 6595 -95
rect 5635 -1465 5755 -170
rect -70 -1510 70 -1500
rect -70 -1530 -60 -1510
rect -10 -1530 70 -1510
rect -70 -1540 70 -1530
rect 6595 -1540 6620 -1500
rect -70 -1595 70 -1555
rect 6595 -1595 6620 -1555
rect 430 -1620 6595 -1610
rect 430 -1640 440 -1620
rect 490 -1640 1240 -1620
rect 1290 -1640 2040 -1620
rect 2090 -1640 2840 -1620
rect 2890 -1640 3640 -1620
rect 3690 -1640 4440 -1620
rect 4490 -1640 5240 -1620
rect 5290 -1640 6595 -1620
rect 430 -1650 6595 -1640
rect 225 -1675 6595 -1665
rect 225 -1695 235 -1675
rect 285 -1695 1035 -1675
rect 1085 -1695 1835 -1675
rect 1885 -1695 2635 -1675
rect 2685 -1695 3435 -1675
rect 3485 -1695 4235 -1675
rect 4285 -1695 5035 -1675
rect 5085 -1695 6595 -1675
rect 225 -1705 6595 -1695
rect -70 -3110 70 -3100
rect -70 -3130 -60 -3110
rect -10 -3130 70 -3110
rect -70 -3140 70 -3130
rect -70 -3195 70 -3155
rect 430 -3220 6490 -3210
rect 430 -3240 440 -3220
rect 490 -3240 1240 -3220
rect 1290 -3240 2040 -3220
rect 2090 -3240 2840 -3220
rect 2890 -3240 3640 -3220
rect 3690 -3240 4440 -3220
rect 4490 -3240 5240 -3220
rect 5290 -3240 6040 -3220
rect 6090 -3240 6490 -3220
rect 430 -3250 6490 -3240
rect 225 -3275 6490 -3265
rect 225 -3295 235 -3275
rect 285 -3295 1035 -3275
rect 1085 -3295 1835 -3275
rect 1885 -3295 2635 -3275
rect 2685 -3295 3435 -3275
rect 3485 -3295 4235 -3275
rect 4285 -3295 5035 -3275
rect 5085 -3295 5835 -3275
rect 5885 -3295 6490 -3275
rect 225 -3305 6490 -3295
rect 5635 -4670 5765 -3375
rect -70 -4715 70 -4705
rect -70 -4735 -60 -4715
rect -10 -4735 70 -4715
rect -70 -4745 70 -4735
rect -70 -4800 70 -4760
rect 430 -4825 5690 -4815
rect 430 -4845 440 -4825
rect 490 -4845 1240 -4825
rect 1290 -4845 2040 -4825
rect 2090 -4845 2840 -4825
rect 2890 -4845 3640 -4825
rect 3690 -4845 4440 -4825
rect 4490 -4845 5240 -4825
rect 5290 -4845 5690 -4825
rect 430 -4855 5690 -4845
rect 225 -4880 5690 -4870
rect 225 -4900 235 -4880
rect 285 -4900 1035 -4880
rect 1085 -4900 1835 -4880
rect 1885 -4900 2635 -4880
rect 2685 -4900 3435 -4880
rect 3485 -4900 4235 -4880
rect 4285 -4900 5035 -4880
rect 5085 -4900 5690 -4880
rect 225 -4910 5690 -4900
rect 4835 -6275 4950 -4980
rect -70 -6320 70 -6310
rect -70 -6340 -60 -6320
rect -10 -6340 70 -6320
rect -70 -6350 70 -6340
rect -70 -6405 70 -6365
rect 430 -6430 6595 -6420
rect 430 -6450 440 -6430
rect 490 -6450 1240 -6430
rect 1290 -6450 2040 -6430
rect 2090 -6450 2840 -6430
rect 2890 -6450 3640 -6430
rect 3690 -6450 4440 -6430
rect 4490 -6450 6595 -6430
rect 430 -6460 6595 -6450
rect 225 -6485 6595 -6475
rect 225 -6505 235 -6485
rect 285 -6505 1035 -6485
rect 1085 -6505 1835 -6485
rect 1885 -6505 2635 -6485
rect 2685 -6505 3435 -6485
rect 3485 -6505 4235 -6485
rect 4285 -6505 6595 -6485
rect 225 -6515 6595 -6505
use dac_unit  dac_unit_0
timestamp 1702614989
transform 1 0 -1115 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_1
timestamp 1702614989
transform 1 0 -315 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_2
timestamp 1702614989
transform 1 0 485 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_3
timestamp 1702614989
transform 1 0 1285 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_4
timestamp 1702614989
transform 1 0 2085 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_5
timestamp 1702614989
transform 1 0 4590 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_6
timestamp 1702614989
transform 1 0 -1115 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_7
timestamp 1702614989
transform 1 0 2085 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_8
timestamp 1702614989
transform 1 0 -315 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_9
timestamp 1702614989
transform 1 0 485 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_10
timestamp 1702614989
transform 1 0 1285 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_11
timestamp 1702614989
transform 1 0 4485 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_12
timestamp 1702614989
transform 1 0 2885 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_13
timestamp 1702614989
transform 1 0 -1115 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_14
timestamp 1702614989
transform 1 0 3685 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_15
timestamp 1702614989
transform 1 0 -315 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_16
timestamp 1702614989
transform 1 0 485 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_17
timestamp 1702614989
transform 1 0 1285 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_18
timestamp 1702614989
transform 1 0 2085 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_19
timestamp 1702614989
transform 1 0 2885 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_20
timestamp 1702614989
transform 1 0 3685 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_21
timestamp 1702614989
transform 1 0 -1115 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_22
timestamp 1702614989
transform 1 0 -315 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_23
timestamp 1702614989
transform 1 0 485 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_24
timestamp 1702614989
transform 1 0 1285 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_25
timestamp 1702614989
transform 1 0 2885 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_26
timestamp 1702614989
transform 1 0 -1115 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_27
timestamp 1702614989
transform 1 0 3685 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_28
timestamp 1702614989
transform 1 0 2085 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_29
timestamp 1702614989
transform 1 0 2885 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_30
timestamp 1702614989
transform 1 0 2885 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_31
timestamp 1702614989
transform 1 0 2085 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_32
timestamp 1702614989
transform 1 0 1285 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_33
timestamp 1702614989
transform 1 0 485 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_34
timestamp 1702614989
transform 1 0 -315 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_35
timestamp 1702614989
transform 1 0 3790 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_36
timestamp 1702614989
transform 1 0 3790 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_37
timestamp 1702614989
transform 1 0 4590 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_38
timestamp 1702614989
transform 1 0 4590 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_40
timestamp 1702614989
transform 1 0 4590 0 1 -50
box 1115 55 2005 1520
<< end >>
