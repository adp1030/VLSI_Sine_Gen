magic
tech sky130A
timestamp 1702769090
<< nwell >>
rect -85 1220 60 1430
rect 0 135 60 1220
rect 5245 105 5350 1460
rect 6155 105 6260 1460
rect -90 -380 65 -170
rect 0 -1255 65 -380
rect -15 -1465 65 -1255
rect 6125 -1495 6230 -140
rect -90 -1980 65 -1770
rect -15 -3065 65 -1980
rect -90 -3580 65 -3370
rect 0 -4460 65 -3580
rect -15 -4670 65 -4460
rect 6120 -4700 6250 -3345
rect 0 -4975 65 -4950
rect -90 -5185 65 -4975
rect 0 -5940 65 -5185
rect -35 -5965 65 -5940
rect -85 -6140 65 -5965
rect -150 -6150 65 -6140
rect -175 -6205 65 -6150
rect -150 -6210 65 -6205
rect -70 -6255 65 -6210
rect -75 -6275 65 -6255
rect 5240 -4980 5345 -4950
rect 6145 -4980 6250 -4950
rect 5240 -6275 5350 -4980
rect 6145 -6275 6255 -4980
rect -75 -6305 60 -6275
rect 5240 -6305 5345 -6275
rect 6145 -6305 6250 -6275
<< poly >>
rect 6455 1575 6505 1585
rect -15 1560 6505 1575
rect -15 -25 0 1560
rect 270 1430 320 1560
rect 370 1520 420 1530
rect 370 1500 380 1520
rect 410 1500 420 1520
rect 370 1430 420 1500
rect 1150 1430 1200 1560
rect 1250 1520 1300 1530
rect 1250 1500 1260 1520
rect 1290 1500 1300 1520
rect 1250 1435 1300 1500
rect 2030 1430 2080 1560
rect 2130 1520 2180 1530
rect 2130 1500 2140 1520
rect 2170 1500 2180 1520
rect 2130 1435 2180 1500
rect 2910 1430 2960 1560
rect 3010 1520 3060 1530
rect 3010 1500 3020 1520
rect 3050 1500 3060 1520
rect 3010 1435 3060 1500
rect 3790 1430 3840 1560
rect 3890 1520 3940 1530
rect 3890 1500 3900 1520
rect 3930 1500 3940 1520
rect 3890 1435 3940 1500
rect 4670 1430 4720 1560
rect 4770 1520 4820 1530
rect 4770 1500 4780 1520
rect 4810 1500 4820 1520
rect 4770 1435 4820 1500
rect 5575 1430 5625 1560
rect 5675 1520 5725 1530
rect 5675 1500 5685 1520
rect 5715 1500 5725 1520
rect 5675 1435 5725 1500
rect 6455 1430 6505 1560
rect 6555 1530 6605 1585
rect 6555 1520 7155 1530
rect 6555 1500 6565 1520
rect 6595 1500 7155 1520
rect 6555 1435 6605 1500
rect -15 -40 6505 -25
rect -15 -1625 0 -40
rect 270 -165 320 -40
rect 1070 -75 1120 -65
rect 1070 -80 1080 -75
rect 370 -95 1080 -80
rect 1110 -95 1120 -75
rect 370 -100 1120 -95
rect 370 -165 420 -100
rect 1070 -105 1120 -100
rect 1150 -165 1200 -40
rect 1250 -75 1300 -65
rect 1250 -95 1260 -75
rect 1290 -80 1300 -75
rect 1950 -75 2000 -65
rect 1950 -80 1960 -75
rect 1290 -95 1960 -80
rect 1990 -95 2000 -75
rect 1250 -100 2000 -95
rect 1250 -165 1300 -100
rect 1950 -105 2000 -100
rect 2030 -165 2080 -40
rect 2130 -75 2180 -65
rect 2130 -95 2140 -75
rect 2170 -80 2180 -75
rect 2830 -75 2880 -65
rect 2830 -80 2840 -75
rect 2170 -95 2840 -80
rect 2870 -95 2880 -75
rect 2130 -100 2880 -95
rect 2130 -165 2180 -100
rect 2830 -105 2880 -100
rect 2910 -165 2960 -40
rect 3010 -75 3060 -65
rect 3010 -95 3020 -75
rect 3050 -80 3060 -75
rect 3710 -75 3760 -65
rect 3710 -80 3720 -75
rect 3050 -95 3720 -80
rect 3750 -95 3760 -75
rect 3010 -100 3760 -95
rect 3010 -165 3060 -100
rect 3710 -105 3760 -100
rect 3790 -165 3840 -40
rect 3890 -75 3940 -65
rect 3890 -95 3900 -75
rect 3930 -80 3940 -75
rect 4590 -75 4640 -65
rect 4590 -80 4600 -75
rect 3930 -95 4600 -80
rect 4630 -95 4640 -75
rect 3890 -100 4640 -95
rect 3890 -165 3940 -100
rect 4590 -105 4640 -100
rect 4670 -165 4720 -40
rect 4770 -75 4820 -65
rect 4770 -95 4780 -75
rect 4810 -80 4820 -75
rect 5470 -75 5520 -65
rect 5470 -80 5480 -75
rect 4810 -95 5480 -80
rect 5510 -95 5520 -75
rect 4770 -100 5520 -95
rect 4770 -165 4820 -100
rect 5470 -105 5520 -100
rect 5550 -165 5600 -40
rect 5650 -75 5700 -65
rect 5650 -95 5660 -75
rect 5690 -80 5700 -75
rect 6375 -75 6425 -65
rect 6375 -80 6385 -75
rect 5690 -95 6385 -80
rect 6415 -95 6425 -75
rect 5650 -100 6425 -95
rect 5650 -165 5700 -100
rect 6375 -105 6425 -100
rect 6455 -165 6505 -40
rect 6555 -75 6605 -65
rect 6555 -95 6565 -75
rect 6595 -80 6605 -75
rect 7120 -80 7155 1500
rect 6595 -95 7155 -80
rect 6555 -100 7155 -95
rect 6555 -165 6605 -100
rect -15 -1640 6480 -1625
rect -15 -3225 0 -1640
rect 270 -1765 320 -1640
rect 370 -1680 420 -1665
rect 1070 -1675 1120 -1665
rect 1070 -1680 1080 -1675
rect 370 -1695 1080 -1680
rect 1110 -1695 1120 -1675
rect 370 -1700 1120 -1695
rect 370 -1765 420 -1700
rect 1070 -1705 1120 -1700
rect 1150 -1765 1200 -1640
rect 1250 -1675 1300 -1665
rect 1250 -1695 1260 -1675
rect 1290 -1680 1300 -1675
rect 1950 -1675 2000 -1665
rect 1950 -1680 1960 -1675
rect 1290 -1695 1960 -1680
rect 1990 -1695 2000 -1675
rect 1250 -1700 2000 -1695
rect 1250 -1765 1300 -1700
rect 1950 -1705 2000 -1700
rect 2030 -1765 2080 -1640
rect 2130 -1675 2180 -1665
rect 2130 -1695 2140 -1675
rect 2170 -1680 2180 -1675
rect 2830 -1675 2880 -1665
rect 2830 -1680 2840 -1675
rect 2170 -1695 2840 -1680
rect 2870 -1695 2880 -1675
rect 2130 -1700 2880 -1695
rect 2130 -1770 2180 -1700
rect 2830 -1705 2880 -1700
rect 2910 -1765 2960 -1640
rect 3010 -1675 3060 -1665
rect 3010 -1695 3020 -1675
rect 3050 -1680 3060 -1675
rect 3710 -1675 3760 -1665
rect 3710 -1680 3720 -1675
rect 3050 -1695 3720 -1680
rect 3750 -1695 3760 -1675
rect 3010 -1700 3760 -1695
rect 3010 -1765 3060 -1700
rect 3710 -1705 3760 -1700
rect 3790 -1765 3840 -1640
rect 3890 -1675 3940 -1665
rect 3890 -1695 3900 -1675
rect 3930 -1680 3940 -1675
rect 4590 -1675 4640 -1665
rect 4590 -1680 4600 -1675
rect 3930 -1695 4600 -1680
rect 4630 -1695 4640 -1675
rect 3890 -1700 4640 -1695
rect 3890 -1765 3940 -1700
rect 4590 -1705 4640 -1700
rect 4670 -1765 4720 -1640
rect 4770 -1675 4820 -1665
rect 4770 -1695 4780 -1675
rect 4810 -1680 4820 -1675
rect 5470 -1675 5520 -1665
rect 5470 -1680 5480 -1675
rect 4810 -1695 5480 -1680
rect 5510 -1695 5520 -1675
rect 4770 -1700 5520 -1695
rect 4770 -1765 4820 -1700
rect 5470 -1705 5520 -1700
rect 5550 -1765 5600 -1640
rect 5650 -1675 5700 -1665
rect 5650 -1695 5660 -1675
rect 5690 -1680 5700 -1675
rect 6350 -1675 6400 -1665
rect 6350 -1680 6360 -1675
rect 5690 -1695 6360 -1680
rect 6390 -1695 6400 -1675
rect 5650 -1700 6400 -1695
rect 5650 -1765 5700 -1700
rect 6350 -1705 6400 -1700
rect 6430 -1765 6480 -1640
rect 6530 -1675 6580 -1665
rect 6530 -1695 6540 -1675
rect 6570 -1680 6580 -1675
rect 7120 -1680 7155 -100
rect 6570 -1695 7155 -1680
rect 6530 -1700 7155 -1695
rect 6530 -1765 6580 -1700
rect -15 -3240 6505 -3225
rect -15 -4830 0 -3240
rect 270 -3370 320 -3240
rect 370 -3280 420 -3265
rect 1070 -3275 1120 -3265
rect 1070 -3280 1080 -3275
rect 370 -3295 1080 -3280
rect 1110 -3295 1120 -3275
rect 370 -3300 1120 -3295
rect 370 -3370 420 -3300
rect 1070 -3305 1120 -3300
rect 1150 -3370 1200 -3240
rect 1250 -3275 1300 -3265
rect 1250 -3295 1260 -3275
rect 1290 -3280 1300 -3275
rect 1950 -3275 2000 -3265
rect 1950 -3280 1960 -3275
rect 1290 -3295 1960 -3280
rect 1990 -3295 2000 -3275
rect 1250 -3300 2000 -3295
rect 1250 -3370 1300 -3300
rect 1950 -3305 2000 -3300
rect 2030 -3375 2080 -3240
rect 2130 -3275 2180 -3265
rect 2130 -3295 2140 -3275
rect 2170 -3280 2180 -3275
rect 2830 -3275 2880 -3265
rect 2830 -3280 2840 -3275
rect 2170 -3295 2840 -3280
rect 2870 -3295 2880 -3275
rect 2130 -3300 2880 -3295
rect 2130 -3370 2180 -3300
rect 2830 -3305 2880 -3300
rect 2910 -3370 2960 -3240
rect 3010 -3275 3060 -3265
rect 3010 -3295 3020 -3275
rect 3050 -3280 3060 -3275
rect 3710 -3275 3760 -3265
rect 3710 -3280 3720 -3275
rect 3050 -3295 3720 -3280
rect 3750 -3295 3760 -3275
rect 3010 -3300 3760 -3295
rect 3010 -3370 3060 -3300
rect 3710 -3305 3760 -3300
rect 3790 -3370 3840 -3240
rect 3890 -3275 3940 -3265
rect 3890 -3295 3900 -3275
rect 3930 -3280 3940 -3275
rect 4590 -3275 4640 -3265
rect 4590 -3280 4600 -3275
rect 3930 -3295 4600 -3280
rect 4630 -3295 4640 -3275
rect 3890 -3300 4640 -3295
rect 3890 -3370 3940 -3300
rect 4590 -3305 4640 -3300
rect 4670 -3370 4720 -3240
rect 4770 -3275 4820 -3265
rect 4770 -3295 4780 -3275
rect 4810 -3280 4820 -3275
rect 5470 -3275 5520 -3265
rect 5470 -3280 5480 -3275
rect 4810 -3295 5480 -3280
rect 5510 -3295 5520 -3275
rect 4770 -3300 5520 -3295
rect 4770 -3370 4820 -3300
rect 5470 -3305 5520 -3300
rect 5550 -3370 5600 -3240
rect 5650 -3275 5700 -3265
rect 5650 -3295 5660 -3275
rect 5690 -3280 5700 -3275
rect 6375 -3275 6425 -3265
rect 6375 -3280 6385 -3275
rect 5690 -3295 6385 -3280
rect 6415 -3295 6425 -3275
rect 5650 -3300 6425 -3295
rect 5650 -3370 5700 -3300
rect 6375 -3305 6425 -3300
rect 6455 -3370 6505 -3240
rect 6555 -3275 6605 -3265
rect 6555 -3295 6565 -3275
rect 6595 -3280 6605 -3275
rect 7120 -3280 7155 -1700
rect 6595 -3295 7155 -3280
rect 6555 -3300 7155 -3295
rect 6555 -3370 6605 -3300
rect -15 -4845 6505 -4830
rect 270 -4975 320 -4845
rect 370 -4885 420 -4870
rect 1070 -4880 1120 -4870
rect 1070 -4885 1080 -4880
rect 370 -4900 1080 -4885
rect 1110 -4900 1120 -4880
rect 370 -4905 1120 -4900
rect 370 -4975 420 -4905
rect 1070 -4910 1120 -4905
rect 1150 -4975 1200 -4845
rect 1250 -4880 1300 -4870
rect 1250 -4900 1260 -4880
rect 1290 -4885 1300 -4880
rect 1950 -4880 2000 -4870
rect 1950 -4885 1960 -4880
rect 1290 -4900 1960 -4885
rect 1990 -4900 2000 -4880
rect 1250 -4905 2000 -4900
rect 1250 -4975 1300 -4905
rect 1950 -4910 2000 -4905
rect 2030 -4975 2080 -4845
rect 2130 -4880 2180 -4870
rect 2130 -4900 2140 -4880
rect 2170 -4885 2180 -4880
rect 2830 -4880 2880 -4870
rect 2830 -4885 2840 -4880
rect 2170 -4900 2840 -4885
rect 2870 -4900 2880 -4880
rect 2130 -4905 2880 -4900
rect 2130 -4975 2180 -4905
rect 2830 -4910 2880 -4905
rect 2910 -4975 2960 -4845
rect 3010 -4880 3060 -4870
rect 3010 -4900 3020 -4880
rect 3050 -4885 3060 -4880
rect 3710 -4880 3760 -4870
rect 3710 -4885 3720 -4880
rect 3050 -4900 3720 -4885
rect 3750 -4900 3760 -4880
rect 3010 -4905 3760 -4900
rect 3010 -4975 3060 -4905
rect 3710 -4910 3760 -4905
rect 3790 -4975 3840 -4845
rect 3890 -4880 3940 -4870
rect 3890 -4900 3900 -4880
rect 3930 -4885 3940 -4880
rect 4590 -4880 4640 -4870
rect 4590 -4885 4600 -4880
rect 3930 -4900 4600 -4885
rect 4630 -4900 4640 -4880
rect 3890 -4905 4640 -4900
rect 3890 -4975 3940 -4905
rect 4590 -4910 4640 -4905
rect 4670 -4975 4720 -4845
rect 4770 -4880 4820 -4870
rect 4770 -4900 4780 -4880
rect 4810 -4885 4820 -4880
rect 5495 -4880 5545 -4870
rect 5495 -4885 5505 -4880
rect 4810 -4900 5505 -4885
rect 5535 -4900 5545 -4880
rect 4770 -4905 5545 -4900
rect 4770 -4975 4820 -4905
rect 5495 -4910 5545 -4905
rect 5575 -4975 5625 -4845
rect 5675 -4880 5725 -4870
rect 5675 -4900 5685 -4880
rect 5715 -4885 5725 -4880
rect 6375 -4880 6425 -4870
rect 6375 -4885 6385 -4880
rect 5715 -4900 6385 -4885
rect 6415 -4900 6425 -4880
rect 5675 -4905 6425 -4900
rect 5675 -4975 5725 -4905
rect 6375 -4910 6425 -4905
rect 6455 -4975 6505 -4845
rect 6555 -4880 6605 -4870
rect 6555 -4900 6565 -4880
rect 6595 -4885 6605 -4880
rect 7120 -4885 7155 -3300
rect 6595 -4900 7155 -4885
rect 6555 -4905 7155 -4900
rect 6555 -4975 6605 -4905
rect -365 -5875 -325 -5865
rect -365 -5895 -355 -5875
rect -335 -5895 -325 -5875
rect -365 -6055 -325 -5895
<< polycont >>
rect 380 1500 410 1520
rect 1260 1500 1290 1520
rect 2140 1500 2170 1520
rect 3020 1500 3050 1520
rect 3900 1500 3930 1520
rect 4780 1500 4810 1520
rect 5685 1500 5715 1520
rect 6565 1500 6595 1520
rect 1080 -95 1110 -75
rect 1260 -95 1290 -75
rect 1960 -95 1990 -75
rect 2140 -95 2170 -75
rect 2840 -95 2870 -75
rect 3020 -95 3050 -75
rect 3720 -95 3750 -75
rect 3900 -95 3930 -75
rect 4600 -95 4630 -75
rect 4780 -95 4810 -75
rect 5480 -95 5510 -75
rect 5660 -95 5690 -75
rect 6385 -95 6415 -75
rect 6565 -95 6595 -75
rect 1080 -1695 1110 -1675
rect 1260 -1695 1290 -1675
rect 1960 -1695 1990 -1675
rect 2140 -1695 2170 -1675
rect 2840 -1695 2870 -1675
rect 3020 -1695 3050 -1675
rect 3720 -1695 3750 -1675
rect 3900 -1695 3930 -1675
rect 4600 -1695 4630 -1675
rect 4780 -1695 4810 -1675
rect 5480 -1695 5510 -1675
rect 5660 -1695 5690 -1675
rect 6360 -1695 6390 -1675
rect 6540 -1695 6570 -1675
rect 1080 -3295 1110 -3275
rect 1260 -3295 1290 -3275
rect 1960 -3295 1990 -3275
rect 2140 -3295 2170 -3275
rect 2840 -3295 2870 -3275
rect 3020 -3295 3050 -3275
rect 3720 -3295 3750 -3275
rect 3900 -3295 3930 -3275
rect 4600 -3295 4630 -3275
rect 4780 -3295 4810 -3275
rect 5480 -3295 5510 -3275
rect 5660 -3295 5690 -3275
rect 6385 -3295 6415 -3275
rect 6565 -3295 6595 -3275
rect 1080 -4900 1110 -4880
rect 1260 -4900 1290 -4880
rect 1960 -4900 1990 -4880
rect 2140 -4900 2170 -4880
rect 2840 -4900 2870 -4880
rect 3020 -4900 3050 -4880
rect 3720 -4900 3750 -4880
rect 3900 -4900 3930 -4880
rect 4600 -4900 4630 -4880
rect 4780 -4900 4810 -4880
rect 5505 -4900 5535 -4880
rect 5685 -4900 5715 -4880
rect 6385 -4900 6415 -4880
rect 6565 -4900 6595 -4880
rect -355 -5895 -335 -5875
<< locali >>
rect -415 1580 80 1590
rect -415 1560 20 1580
rect 70 1560 80 1580
rect -415 1550 80 1560
rect -405 1240 -385 1550
rect -345 1520 80 1530
rect -345 1500 20 1520
rect 70 1500 80 1520
rect -345 1490 80 1500
rect 370 1520 6605 1530
rect 370 1500 380 1520
rect 410 1500 1260 1520
rect 1290 1500 2140 1520
rect 2170 1500 3020 1520
rect 3050 1500 3900 1520
rect 3930 1500 4780 1520
rect 4810 1500 5685 1520
rect 5715 1500 6565 1520
rect 6595 1500 6605 1520
rect 370 1495 6605 1500
rect 370 1490 420 1495
rect 1250 1490 1300 1495
rect 2130 1490 2180 1495
rect 3010 1490 3060 1495
rect 3890 1490 3940 1495
rect 4770 1490 4820 1495
rect 5675 1490 5725 1495
rect 6555 1490 6605 1495
rect -345 1405 -325 1490
rect -405 1220 -325 1240
rect 7145 175 7185 185
rect 7145 125 7155 175
rect 7175 125 7185 175
rect -415 90 80 100
rect -415 70 20 90
rect 70 70 80 90
rect -415 60 80 70
rect -405 -360 -385 60
rect -345 30 80 40
rect -345 10 20 30
rect 70 10 80 30
rect -345 0 80 10
rect -345 -195 -325 0
rect 225 -65 260 45
rect 430 -10 460 45
rect 430 -20 500 -10
rect 430 -40 440 -20
rect 490 -40 500 -20
rect 430 -50 500 -40
rect 1000 -15 1140 20
rect 1310 -10 1340 45
rect 1985 20 2020 45
rect 1000 -65 1035 -15
rect 1310 -20 1380 -10
rect 1310 -40 1320 -20
rect 1370 -40 1380 -20
rect 1310 -50 1380 -40
rect 1880 -15 2020 20
rect 2190 -10 2220 45
rect 2865 20 2900 45
rect 1880 -65 1915 -15
rect 2190 -20 2260 -10
rect 2190 -40 2200 -20
rect 2250 -40 2260 -20
rect 2190 -50 2260 -40
rect 2760 -15 2900 20
rect 3070 -10 3100 45
rect 3745 20 3780 45
rect 2760 -65 2795 -15
rect 3070 -20 3140 -10
rect 3070 -40 3080 -20
rect 3130 -40 3140 -20
rect 3070 -50 3140 -40
rect 3640 -15 3780 20
rect 3950 -10 3980 45
rect 4625 20 4660 45
rect 3640 -65 3675 -15
rect 3950 -20 4020 -10
rect 3950 -40 3960 -20
rect 4010 -40 4020 -20
rect 3950 -50 4020 -40
rect 4520 -15 4660 20
rect 4830 -10 4860 45
rect 5535 20 5565 45
rect 4520 -65 4555 -15
rect 4830 -20 4900 -10
rect 4830 -40 4840 -20
rect 4890 -40 4900 -20
rect 4830 -50 4900 -40
rect 5405 -15 5565 20
rect 5735 -10 5765 45
rect 6435 20 6445 45
rect 5735 -15 5785 -10
rect 5405 -65 5440 -15
rect 5715 -20 5785 -15
rect 5715 -40 5725 -20
rect 5775 -40 5785 -20
rect 5715 -50 5785 -40
rect 6305 -15 6445 20
rect 6615 -10 6645 50
rect 7145 45 7185 125
rect 7115 40 7185 45
rect 7115 20 7125 40
rect 7175 20 7185 40
rect 7115 10 7185 20
rect 6305 -65 6340 -15
rect 6615 -20 6685 -10
rect 6615 -40 6625 -20
rect 6675 -40 6685 -20
rect 6615 -50 6685 -40
rect 7060 -20 7350 -10
rect 7060 -40 7070 -20
rect 7120 -40 7290 -20
rect 7340 -40 7350 -20
rect 7060 -50 7350 -40
rect 225 -75 295 -65
rect 225 -95 235 -75
rect 285 -95 295 -75
rect 225 -105 295 -95
rect 965 -75 1035 -65
rect 965 -95 975 -75
rect 1025 -95 1035 -75
rect 965 -105 1035 -95
rect 1070 -75 1300 -65
rect 1070 -95 1080 -75
rect 1110 -95 1260 -75
rect 1290 -95 1300 -75
rect 1070 -105 1300 -95
rect 1845 -75 1915 -65
rect 1845 -95 1855 -75
rect 1905 -95 1915 -75
rect 1845 -105 1915 -95
rect 1950 -75 2180 -65
rect 1950 -95 1960 -75
rect 1990 -95 2140 -75
rect 2170 -95 2180 -75
rect 1950 -105 2180 -95
rect 2725 -75 2795 -65
rect 2725 -95 2735 -75
rect 2785 -95 2795 -75
rect 2725 -105 2795 -95
rect 2830 -75 3060 -65
rect 2830 -95 2840 -75
rect 2870 -95 3020 -75
rect 3050 -95 3060 -75
rect 2830 -105 3060 -95
rect 3605 -75 3675 -65
rect 3605 -95 3615 -75
rect 3665 -95 3675 -75
rect 3605 -105 3675 -95
rect 3710 -75 3940 -65
rect 3710 -95 3720 -75
rect 3750 -95 3900 -75
rect 3930 -95 3940 -75
rect 3710 -105 3940 -95
rect 4485 -75 4555 -65
rect 4485 -95 4495 -75
rect 4545 -95 4555 -75
rect 4485 -105 4555 -95
rect 4590 -75 4820 -65
rect 4590 -95 4600 -75
rect 4630 -95 4780 -75
rect 4810 -95 4820 -75
rect 4590 -105 4820 -95
rect 5370 -75 5440 -65
rect 5370 -95 5380 -75
rect 5430 -95 5440 -75
rect 5370 -105 5440 -95
rect 5470 -75 5700 -65
rect 5470 -95 5480 -75
rect 5510 -95 5660 -75
rect 5690 -95 5700 -75
rect 5470 -105 5700 -95
rect 6270 -75 6340 -65
rect 6270 -95 6280 -75
rect 6330 -95 6340 -75
rect 6270 -105 6340 -95
rect 6375 -75 6605 -65
rect 6375 -95 6385 -75
rect 6415 -95 6565 -75
rect 6595 -95 6605 -75
rect 6375 -105 6605 -95
rect 7090 -85 7130 -75
rect 7090 -135 7100 -85
rect 7120 -105 7130 -85
rect 7120 -115 7295 -105
rect 7120 -135 7265 -115
rect 7090 -145 7265 -135
rect 7255 -165 7265 -145
rect 7285 -165 7295 -115
rect 7255 -175 7295 -165
rect -405 -380 -325 -360
rect 7200 -1450 7240 -1440
rect 7200 -1475 7210 -1450
rect 7090 -1500 7210 -1475
rect 7230 -1500 7240 -1450
rect -415 -1510 80 -1500
rect -415 -1530 20 -1510
rect 70 -1530 80 -1510
rect -415 -1540 80 -1530
rect 7050 -1510 7240 -1500
rect 7050 -1530 7065 -1510
rect 7115 -1530 7130 -1510
rect 7050 -1540 7130 -1530
rect 7255 -1535 7295 -1525
rect -405 -1960 -385 -1540
rect -345 -1570 80 -1560
rect -345 -1590 20 -1570
rect 70 -1590 80 -1570
rect -345 -1600 80 -1590
rect -345 -1795 -325 -1600
rect 225 -1665 260 -1555
rect 430 -1610 460 -1555
rect 430 -1620 500 -1610
rect 430 -1640 440 -1620
rect 490 -1640 500 -1620
rect 430 -1650 500 -1640
rect 1000 -1615 1140 -1580
rect 1310 -1610 1340 -1555
rect 1000 -1665 1035 -1615
rect 1310 -1620 1380 -1610
rect 1310 -1640 1320 -1620
rect 1370 -1640 1380 -1620
rect 1310 -1650 1380 -1640
rect 1880 -1615 2020 -1580
rect 2190 -1610 2220 -1555
rect 1880 -1665 1915 -1615
rect 2190 -1620 2260 -1610
rect 2190 -1640 2200 -1620
rect 2250 -1640 2260 -1620
rect 2190 -1650 2260 -1640
rect 2760 -1615 2900 -1580
rect 3070 -1610 3100 -1555
rect 2760 -1665 2795 -1615
rect 3070 -1620 3140 -1610
rect 3070 -1640 3080 -1620
rect 3130 -1640 3140 -1620
rect 3070 -1650 3140 -1640
rect 3640 -1615 3780 -1580
rect 3950 -1610 3980 -1555
rect 3640 -1665 3675 -1615
rect 3950 -1620 4020 -1610
rect 3950 -1640 3960 -1620
rect 4010 -1640 4020 -1620
rect 3950 -1650 4020 -1640
rect 4520 -1615 4660 -1580
rect 4830 -1610 4860 -1555
rect 5535 -1580 5540 -1550
rect 4520 -1665 4555 -1615
rect 4835 -1620 4905 -1610
rect 4835 -1640 4845 -1620
rect 4895 -1640 4905 -1620
rect 4835 -1650 4905 -1640
rect 5410 -1615 5540 -1580
rect 5710 -1610 5740 -1555
rect 6420 -1580 6445 -1555
rect 5410 -1665 5445 -1615
rect 5715 -1620 5785 -1610
rect 5715 -1640 5725 -1620
rect 5775 -1640 5785 -1620
rect 5715 -1650 5785 -1640
rect 6270 -1615 6445 -1580
rect 6615 -1610 6645 -1545
rect 7255 -1585 7265 -1535
rect 7285 -1585 7295 -1535
rect 6270 -1665 6305 -1615
rect 6595 -1620 6665 -1610
rect 6595 -1640 6605 -1620
rect 6655 -1640 6665 -1620
rect 6595 -1650 6665 -1640
rect 225 -1675 295 -1665
rect 225 -1695 235 -1675
rect 285 -1695 295 -1675
rect 225 -1705 295 -1695
rect 965 -1675 1035 -1665
rect 965 -1695 975 -1675
rect 1025 -1695 1035 -1675
rect 965 -1705 1035 -1695
rect 1070 -1675 1300 -1665
rect 1070 -1695 1080 -1675
rect 1110 -1695 1260 -1675
rect 1290 -1695 1300 -1675
rect 1070 -1705 1300 -1695
rect 1845 -1675 1915 -1665
rect 1845 -1695 1855 -1675
rect 1905 -1695 1915 -1675
rect 1845 -1705 1915 -1695
rect 1950 -1675 2180 -1665
rect 1950 -1695 1960 -1675
rect 1990 -1695 2140 -1675
rect 2170 -1695 2180 -1675
rect 1950 -1705 2180 -1695
rect 2725 -1675 2795 -1665
rect 2725 -1695 2735 -1675
rect 2785 -1695 2795 -1675
rect 2725 -1705 2795 -1695
rect 2830 -1675 3060 -1665
rect 2830 -1695 2840 -1675
rect 2870 -1695 3020 -1675
rect 3050 -1695 3060 -1675
rect 2830 -1705 3060 -1695
rect 3605 -1675 3675 -1665
rect 3605 -1695 3615 -1675
rect 3665 -1695 3675 -1675
rect 3605 -1705 3675 -1695
rect 3710 -1675 3940 -1665
rect 3710 -1695 3720 -1675
rect 3750 -1695 3900 -1675
rect 3930 -1695 3940 -1675
rect 3710 -1705 3940 -1695
rect 4485 -1675 4555 -1665
rect 4485 -1695 4495 -1675
rect 4545 -1695 4555 -1675
rect 4485 -1705 4555 -1695
rect 4590 -1675 4820 -1665
rect 4590 -1695 4600 -1675
rect 4630 -1695 4780 -1675
rect 4810 -1695 4820 -1675
rect 4590 -1705 4820 -1695
rect 5375 -1675 5445 -1665
rect 5375 -1695 5385 -1675
rect 5435 -1695 5445 -1675
rect 5375 -1705 5445 -1695
rect 5470 -1675 5700 -1665
rect 5470 -1695 5480 -1675
rect 5510 -1695 5660 -1675
rect 5690 -1695 5700 -1675
rect 5470 -1705 5700 -1695
rect 6235 -1675 6305 -1665
rect 6235 -1695 6245 -1675
rect 6295 -1695 6305 -1675
rect 6235 -1705 6305 -1695
rect 6350 -1675 6580 -1665
rect 6350 -1695 6360 -1675
rect 6390 -1695 6540 -1675
rect 6570 -1695 6580 -1675
rect 6350 -1705 6580 -1695
rect 7255 -1675 7295 -1585
rect 7255 -1725 7265 -1675
rect 7285 -1725 7295 -1675
rect 7255 -1740 7295 -1725
rect -405 -1980 -325 -1960
rect -415 -3110 80 -3100
rect -415 -3130 20 -3110
rect 70 -3130 80 -3110
rect -415 -3140 80 -3130
rect 7255 -3135 7295 -3125
rect -405 -3560 -385 -3140
rect -345 -3170 80 -3160
rect -345 -3190 20 -3170
rect 70 -3190 80 -3170
rect -345 -3200 80 -3190
rect -345 -3395 -325 -3200
rect 225 -3265 260 -3155
rect 430 -3210 460 -3155
rect 430 -3220 500 -3210
rect 430 -3240 440 -3220
rect 490 -3240 500 -3220
rect 430 -3250 500 -3240
rect 1000 -3215 1140 -3180
rect 1310 -3210 1340 -3155
rect 1000 -3265 1035 -3215
rect 1310 -3220 1380 -3210
rect 1310 -3240 1320 -3220
rect 1370 -3240 1380 -3220
rect 1310 -3250 1380 -3240
rect 1880 -3215 2020 -3180
rect 2190 -3210 2220 -3155
rect 1880 -3265 1915 -3215
rect 2190 -3220 2260 -3210
rect 2190 -3240 2200 -3220
rect 2250 -3240 2260 -3220
rect 2190 -3250 2260 -3240
rect 2760 -3215 2900 -3180
rect 3070 -3210 3100 -3155
rect 2760 -3265 2795 -3215
rect 3070 -3220 3140 -3210
rect 3070 -3240 3080 -3220
rect 3130 -3240 3140 -3220
rect 3070 -3250 3140 -3240
rect 3640 -3215 3780 -3180
rect 3950 -3210 3980 -3155
rect 4655 -3180 4660 -3160
rect 3640 -3265 3675 -3215
rect 3950 -3220 4020 -3210
rect 3950 -3240 3960 -3220
rect 4010 -3240 4020 -3220
rect 3950 -3250 4020 -3240
rect 4520 -3215 4660 -3180
rect 4830 -3210 4860 -3155
rect 5710 -3170 5735 -3155
rect 6615 -3165 6620 -3155
rect 5535 -3180 5540 -3175
rect 4520 -3265 4555 -3215
rect 4830 -3220 4900 -3210
rect 4830 -3240 4840 -3220
rect 4890 -3240 4900 -3220
rect 4830 -3250 4900 -3240
rect 5410 -3215 5540 -3180
rect 5710 -3210 5740 -3170
rect 6410 -3190 6420 -3175
rect 6615 -3185 6645 -3165
rect 5410 -3265 5445 -3215
rect 5710 -3220 5780 -3210
rect 5710 -3240 5720 -3220
rect 5770 -3240 5780 -3220
rect 5710 -3250 5780 -3240
rect 6295 -3225 6420 -3190
rect 6590 -3210 6645 -3185
rect 7255 -3185 7265 -3135
rect 7285 -3185 7295 -3135
rect 6615 -3220 6690 -3210
rect 6295 -3265 6330 -3225
rect 6615 -3240 6625 -3220
rect 6675 -3240 6690 -3220
rect 6615 -3250 6690 -3240
rect 225 -3275 295 -3265
rect 225 -3295 235 -3275
rect 285 -3295 295 -3275
rect 225 -3305 295 -3295
rect 965 -3275 1035 -3265
rect 965 -3295 975 -3275
rect 1025 -3295 1035 -3275
rect 965 -3305 1035 -3295
rect 1070 -3275 1300 -3265
rect 1070 -3295 1080 -3275
rect 1110 -3295 1260 -3275
rect 1290 -3295 1300 -3275
rect 1070 -3305 1300 -3295
rect 1845 -3275 1915 -3265
rect 1845 -3295 1855 -3275
rect 1905 -3295 1915 -3275
rect 1845 -3305 1915 -3295
rect 1950 -3275 2180 -3265
rect 1950 -3295 1960 -3275
rect 1990 -3295 2140 -3275
rect 2170 -3295 2180 -3275
rect 1950 -3305 2180 -3295
rect 2725 -3275 2795 -3265
rect 2725 -3295 2735 -3275
rect 2785 -3295 2795 -3275
rect 2725 -3305 2795 -3295
rect 2830 -3275 3060 -3265
rect 2830 -3295 2840 -3275
rect 2870 -3295 3020 -3275
rect 3050 -3295 3060 -3275
rect 2830 -3305 3060 -3295
rect 3605 -3275 3675 -3265
rect 3605 -3295 3615 -3275
rect 3665 -3295 3675 -3275
rect 3605 -3305 3675 -3295
rect 3710 -3275 3940 -3265
rect 3710 -3295 3720 -3275
rect 3750 -3295 3900 -3275
rect 3930 -3295 3940 -3275
rect 3710 -3305 3940 -3295
rect 4485 -3275 4555 -3265
rect 4485 -3295 4495 -3275
rect 4545 -3295 4555 -3275
rect 4485 -3305 4555 -3295
rect 4590 -3275 4820 -3265
rect 4590 -3295 4600 -3275
rect 4630 -3295 4780 -3275
rect 4810 -3295 4820 -3275
rect 4590 -3305 4820 -3295
rect 5375 -3275 5445 -3265
rect 5375 -3295 5385 -3275
rect 5435 -3295 5445 -3275
rect 5375 -3305 5445 -3295
rect 5470 -3275 5700 -3265
rect 5470 -3295 5480 -3275
rect 5510 -3295 5660 -3275
rect 5690 -3295 5700 -3275
rect 5470 -3305 5700 -3295
rect 6245 -3275 6330 -3265
rect 6245 -3295 6260 -3275
rect 6320 -3295 6330 -3275
rect 6245 -3305 6330 -3295
rect 6375 -3270 6425 -3265
rect 6555 -3270 6605 -3265
rect 6375 -3275 6605 -3270
rect 6375 -3295 6385 -3275
rect 6415 -3295 6565 -3275
rect 6595 -3295 6605 -3275
rect 6375 -3305 6605 -3295
rect 7255 -3275 7295 -3185
rect 7255 -3325 7265 -3275
rect 7285 -3325 7295 -3275
rect 7255 -3340 7295 -3325
rect -405 -3580 -325 -3560
rect -415 -4715 80 -4705
rect -415 -4735 20 -4715
rect 70 -4735 80 -4715
rect -415 -4745 80 -4735
rect 7180 -4740 7220 -4730
rect -405 -5165 -385 -4745
rect -345 -4775 85 -4765
rect -345 -4795 25 -4775
rect 75 -4795 85 -4775
rect -345 -4805 85 -4795
rect -345 -5000 -325 -4805
rect 225 -4870 260 -4760
rect 430 -4815 460 -4760
rect 430 -4825 500 -4815
rect 430 -4845 440 -4825
rect 490 -4845 500 -4825
rect 430 -4855 500 -4845
rect 1000 -4820 1140 -4790
rect 1310 -4815 1340 -4760
rect 1000 -4870 1035 -4820
rect 1310 -4825 1380 -4815
rect 1310 -4845 1320 -4825
rect 1370 -4845 1380 -4825
rect 1310 -4855 1380 -4845
rect 1880 -4820 2020 -4790
rect 2190 -4815 2220 -4760
rect 1880 -4870 1915 -4820
rect 2190 -4825 2260 -4815
rect 2190 -4845 2200 -4825
rect 2250 -4845 2260 -4825
rect 2190 -4855 2260 -4845
rect 2760 -4820 2900 -4790
rect 3070 -4815 3100 -4760
rect 2760 -4870 2795 -4820
rect 3070 -4825 3140 -4815
rect 3070 -4845 3080 -4825
rect 3130 -4845 3140 -4825
rect 3070 -4855 3140 -4845
rect 3640 -4820 3780 -4790
rect 3950 -4815 3980 -4760
rect 3640 -4870 3675 -4820
rect 3950 -4825 4020 -4815
rect 3950 -4845 3960 -4825
rect 4010 -4845 4020 -4825
rect 3950 -4855 4020 -4845
rect 4520 -4820 4660 -4790
rect 4830 -4815 4860 -4760
rect 5735 -4765 5740 -4760
rect 4520 -4870 4555 -4820
rect 4830 -4825 4900 -4815
rect 4830 -4845 4840 -4825
rect 4890 -4845 4900 -4825
rect 4830 -4855 4900 -4845
rect 5425 -4825 5540 -4790
rect 5735 -4815 5765 -4765
rect 6385 -4790 6420 -4755
rect 7090 -4770 7160 -4760
rect 5735 -4825 5810 -4815
rect 5425 -4870 5460 -4825
rect 5735 -4845 5745 -4825
rect 5795 -4845 5810 -4825
rect 5735 -4855 5810 -4845
rect 6305 -4820 6420 -4790
rect 6615 -4815 6645 -4775
rect 7090 -4790 7100 -4770
rect 7150 -4790 7160 -4770
rect 7090 -4800 7160 -4790
rect 6305 -4870 6340 -4820
rect 6615 -4825 6685 -4815
rect 6615 -4845 6625 -4825
rect 6675 -4845 6685 -4825
rect 6615 -4855 6685 -4845
rect 225 -4880 295 -4870
rect 225 -4900 235 -4880
rect 285 -4900 295 -4880
rect 225 -4910 295 -4900
rect 965 -4880 1035 -4870
rect 965 -4900 975 -4880
rect 1025 -4900 1035 -4880
rect 965 -4910 1035 -4900
rect 1070 -4880 1300 -4870
rect 1070 -4900 1080 -4880
rect 1110 -4900 1260 -4880
rect 1290 -4900 1300 -4880
rect 1070 -4910 1300 -4900
rect 1845 -4880 1915 -4870
rect 1845 -4900 1855 -4880
rect 1905 -4900 1915 -4880
rect 1845 -4910 1915 -4900
rect 1950 -4880 2180 -4870
rect 1950 -4900 1960 -4880
rect 1990 -4900 2140 -4880
rect 2170 -4900 2180 -4880
rect 1950 -4910 2180 -4900
rect 2725 -4880 2795 -4870
rect 2725 -4900 2735 -4880
rect 2785 -4900 2795 -4880
rect 2725 -4910 2795 -4900
rect 2830 -4880 3060 -4870
rect 2830 -4900 2840 -4880
rect 2870 -4900 3020 -4880
rect 3050 -4900 3060 -4880
rect 2830 -4910 3060 -4900
rect 3605 -4880 3675 -4870
rect 3605 -4900 3615 -4880
rect 3665 -4900 3675 -4880
rect 3605 -4910 3675 -4900
rect 3710 -4880 3940 -4870
rect 3710 -4900 3720 -4880
rect 3750 -4900 3900 -4880
rect 3930 -4900 3940 -4880
rect 3710 -4910 3940 -4900
rect 4485 -4880 4555 -4870
rect 4485 -4900 4495 -4880
rect 4545 -4900 4555 -4880
rect 4485 -4910 4555 -4900
rect 4590 -4880 4820 -4870
rect 4590 -4900 4600 -4880
rect 4630 -4900 4780 -4880
rect 4810 -4900 4820 -4880
rect 4590 -4910 4820 -4900
rect 5390 -4880 5460 -4870
rect 5390 -4900 5400 -4880
rect 5450 -4900 5460 -4880
rect 5390 -4910 5460 -4900
rect 5495 -4875 5545 -4870
rect 5675 -4875 5725 -4870
rect 5495 -4880 5725 -4875
rect 5495 -4900 5505 -4880
rect 5535 -4900 5685 -4880
rect 5715 -4900 5725 -4880
rect 5495 -4910 5725 -4900
rect 6275 -4880 6340 -4870
rect 6275 -4900 6285 -4880
rect 6330 -4900 6340 -4880
rect 6275 -4910 6340 -4900
rect 6375 -4880 6605 -4870
rect 6375 -4900 6385 -4880
rect 6415 -4900 6565 -4880
rect 6595 -4900 6605 -4880
rect 6375 -4910 6605 -4900
rect 7120 -4935 7160 -4800
rect 7120 -4985 7130 -4935
rect 7150 -4985 7160 -4935
rect 7120 -4995 7160 -4985
rect 7180 -4790 7190 -4740
rect 7210 -4790 7220 -4740
rect 7180 -4935 7220 -4790
rect 7180 -4985 7190 -4935
rect 7210 -4985 7220 -4935
rect 7255 -4740 7295 -4730
rect 7255 -4790 7265 -4740
rect 7285 -4790 7295 -4740
rect 7255 -4880 7295 -4790
rect 7255 -4930 7265 -4880
rect 7285 -4930 7295 -4880
rect 7255 -4940 7295 -4930
rect 7180 -4995 7220 -4985
rect -405 -5185 -325 -5165
rect -415 -5875 -325 -5865
rect -415 -5895 -355 -5875
rect -335 -5895 -325 -5875
rect -365 -5905 -325 -5895
rect -405 -5955 -325 -5930
rect -405 -6190 -385 -5955
rect -365 -6150 -330 -6050
rect -365 -6170 40 -6150
rect -405 -6210 -20 -6190
rect -40 -6370 -20 -6210
rect 0 -6310 40 -6170
rect 7120 -6235 7160 -6225
rect 7120 -6285 7130 -6235
rect 7150 -6285 7160 -6235
rect 0 -6320 80 -6310
rect 0 -6340 20 -6320
rect 70 -6340 80 -6320
rect 0 -6350 80 -6340
rect -40 -6380 80 -6370
rect -40 -6400 20 -6380
rect 70 -6400 80 -6380
rect -40 -6410 80 -6400
rect 225 -6475 260 -6365
rect 430 -6420 460 -6365
rect 430 -6430 500 -6420
rect 430 -6450 440 -6430
rect 490 -6450 500 -6430
rect 430 -6460 500 -6450
rect 1105 -6475 1140 -6365
rect 1310 -6420 1340 -6365
rect 1310 -6430 1380 -6420
rect 1310 -6450 1320 -6430
rect 1370 -6450 1380 -6430
rect 1310 -6460 1380 -6450
rect 1985 -6475 2020 -6365
rect 2190 -6420 2220 -6365
rect 2190 -6430 2260 -6420
rect 2190 -6450 2200 -6430
rect 2250 -6450 2260 -6430
rect 2190 -6460 2260 -6450
rect 2865 -6475 2900 -6365
rect 3070 -6420 3100 -6365
rect 3070 -6430 3140 -6420
rect 3070 -6450 3080 -6430
rect 3130 -6450 3140 -6430
rect 3070 -6460 3140 -6450
rect 3745 -6475 3780 -6365
rect 3950 -6420 3980 -6365
rect 3950 -6430 4020 -6420
rect 3950 -6450 3960 -6430
rect 4010 -6450 4020 -6430
rect 3950 -6460 4020 -6450
rect 4625 -6475 4660 -6365
rect 4830 -6420 4860 -6365
rect 4830 -6430 4900 -6420
rect 4830 -6450 4840 -6430
rect 4890 -6450 4900 -6430
rect 4830 -6460 4900 -6450
rect 5530 -6475 5565 -6355
rect 5735 -6420 5765 -6355
rect 6640 -6365 6645 -6355
rect 7120 -6365 7160 -6285
rect 5735 -6430 5805 -6420
rect 5735 -6450 5745 -6430
rect 5795 -6450 5805 -6430
rect 5735 -6460 5805 -6450
rect 6410 -6475 6445 -6365
rect 6615 -6420 6645 -6365
rect 7090 -6375 7160 -6365
rect 7090 -6395 7100 -6375
rect 7150 -6395 7160 -6375
rect 7090 -6405 7160 -6395
rect 6615 -6430 6685 -6420
rect 6615 -6450 6625 -6430
rect 6675 -6450 6685 -6430
rect 6615 -6460 6685 -6450
rect 225 -6485 295 -6475
rect -380 -6525 -145 -6495
rect -75 -6515 80 -6495
rect 225 -6505 235 -6485
rect 285 -6505 295 -6485
rect 225 -6515 295 -6505
rect 1105 -6485 1175 -6475
rect 1105 -6505 1115 -6485
rect 1165 -6505 1175 -6485
rect 1105 -6515 1175 -6505
rect 1985 -6485 2055 -6475
rect 1985 -6505 1995 -6485
rect 2045 -6505 2055 -6485
rect 1985 -6515 2055 -6505
rect 2865 -6485 2935 -6475
rect 2865 -6505 2875 -6485
rect 2925 -6505 2935 -6485
rect 2865 -6515 2935 -6505
rect 3745 -6485 3815 -6475
rect 3745 -6505 3755 -6485
rect 3805 -6505 3815 -6485
rect 3745 -6515 3815 -6505
rect 4625 -6485 4695 -6475
rect 4625 -6505 4635 -6485
rect 4685 -6505 4695 -6485
rect 4625 -6515 4695 -6505
rect 5530 -6485 5600 -6475
rect 5530 -6505 5540 -6485
rect 5590 -6505 5600 -6485
rect 5530 -6515 5600 -6505
rect 6410 -6485 6480 -6475
rect 6410 -6505 6420 -6485
rect 6470 -6505 6480 -6485
rect 6410 -6515 6480 -6505
rect -185 -6585 -145 -6525
rect 0 -6535 80 -6515
rect 7120 -6530 7160 -6405
rect 0 -6555 20 -6535
rect 70 -6555 80 -6535
rect 0 -6565 80 -6555
rect 7090 -6540 7160 -6530
rect 7090 -6560 7100 -6540
rect 7150 -6560 7160 -6540
rect 7090 -6570 7160 -6560
rect 7180 -6345 7220 -6335
rect 7180 -6395 7190 -6345
rect 7210 -6395 7220 -6345
rect 7180 -6565 7220 -6395
rect 7255 -6345 7295 -6335
rect 7255 -6395 7265 -6345
rect 7285 -6395 7295 -6345
rect 7255 -6475 7295 -6395
rect 7255 -6485 7330 -6475
rect 7255 -6505 7270 -6485
rect 7320 -6505 7330 -6485
rect 7255 -6515 7330 -6505
rect -185 -6595 80 -6585
rect -185 -6615 20 -6595
rect 70 -6615 80 -6595
rect -185 -6625 80 -6615
rect 7180 -6615 7190 -6565
rect 7210 -6615 7220 -6565
rect 7180 -6625 7220 -6615
<< viali >>
rect 20 1560 70 1580
rect 20 1500 70 1520
rect 7155 125 7175 175
rect 20 70 70 90
rect 20 10 70 30
rect 440 -40 490 -20
rect 1320 -40 1370 -20
rect 2200 -40 2250 -20
rect 3080 -40 3130 -20
rect 3960 -40 4010 -20
rect 4840 -40 4890 -20
rect 5725 -40 5775 -20
rect 7125 20 7175 40
rect 6625 -40 6675 -20
rect 7070 -40 7120 -20
rect 7290 -40 7340 -20
rect 235 -95 285 -75
rect 975 -95 1025 -75
rect 1855 -95 1905 -75
rect 2735 -95 2785 -75
rect 3615 -95 3665 -75
rect 4495 -95 4545 -75
rect 5380 -95 5430 -75
rect 6280 -95 6330 -75
rect 7100 -135 7120 -85
rect 7265 -165 7285 -115
rect 7210 -1500 7230 -1450
rect 20 -1530 70 -1510
rect 7065 -1530 7115 -1510
rect 20 -1590 70 -1570
rect 440 -1640 490 -1620
rect 1320 -1640 1370 -1620
rect 2200 -1640 2250 -1620
rect 3080 -1640 3130 -1620
rect 3960 -1640 4010 -1620
rect 4845 -1640 4895 -1620
rect 5725 -1640 5775 -1620
rect 7265 -1585 7285 -1535
rect 6605 -1640 6655 -1620
rect 235 -1695 285 -1675
rect 975 -1695 1025 -1675
rect 1855 -1695 1905 -1675
rect 2735 -1695 2785 -1675
rect 3615 -1695 3665 -1675
rect 4495 -1695 4545 -1675
rect 5385 -1695 5435 -1675
rect 6245 -1695 6295 -1675
rect 7265 -1725 7285 -1675
rect 20 -3130 70 -3110
rect 20 -3190 70 -3170
rect 440 -3240 490 -3220
rect 1320 -3240 1370 -3220
rect 2200 -3240 2250 -3220
rect 3080 -3240 3130 -3220
rect 3960 -3240 4010 -3220
rect 4840 -3240 4890 -3220
rect 5720 -3240 5770 -3220
rect 7265 -3185 7285 -3135
rect 6625 -3240 6675 -3220
rect 235 -3295 285 -3275
rect 975 -3295 1025 -3275
rect 1855 -3295 1905 -3275
rect 2735 -3295 2785 -3275
rect 3615 -3295 3665 -3275
rect 4495 -3295 4545 -3275
rect 5385 -3295 5435 -3275
rect 6260 -3295 6320 -3275
rect 7265 -3325 7285 -3275
rect 20 -4735 70 -4715
rect 25 -4795 75 -4775
rect 440 -4845 490 -4825
rect 1320 -4845 1370 -4825
rect 2200 -4845 2250 -4825
rect 3080 -4845 3130 -4825
rect 3960 -4845 4010 -4825
rect 4840 -4845 4890 -4825
rect 5745 -4845 5795 -4825
rect 7100 -4790 7150 -4770
rect 6625 -4845 6675 -4825
rect 235 -4900 285 -4880
rect 975 -4900 1025 -4880
rect 1855 -4900 1905 -4880
rect 2735 -4900 2785 -4880
rect 3615 -4900 3665 -4880
rect 4495 -4900 4545 -4880
rect 5400 -4900 5450 -4880
rect 6285 -4900 6330 -4880
rect 7130 -4985 7150 -4935
rect 7190 -4790 7210 -4740
rect 7190 -4985 7210 -4935
rect 7265 -4790 7285 -4740
rect 7265 -4930 7285 -4880
rect 7130 -6285 7150 -6235
rect 20 -6340 70 -6320
rect 20 -6400 70 -6380
rect 440 -6450 490 -6430
rect 1320 -6450 1370 -6430
rect 2200 -6450 2250 -6430
rect 3080 -6450 3130 -6430
rect 3960 -6450 4010 -6430
rect 4840 -6450 4890 -6430
rect 5745 -6450 5795 -6430
rect 7100 -6395 7150 -6375
rect 6625 -6450 6675 -6430
rect 235 -6505 285 -6485
rect 1115 -6505 1165 -6485
rect 1995 -6505 2045 -6485
rect 2875 -6505 2925 -6485
rect 3755 -6505 3805 -6485
rect 4635 -6505 4685 -6485
rect 5540 -6505 5590 -6485
rect 6420 -6505 6470 -6485
rect 20 -6555 70 -6535
rect 7100 -6560 7150 -6540
rect 7190 -6395 7210 -6345
rect 7265 -6395 7285 -6345
rect 7270 -6505 7320 -6485
rect 20 -6615 70 -6595
rect 7190 -6615 7210 -6565
<< metal1 >>
rect 0 1585 80 1590
rect 0 1580 7240 1585
rect 0 1560 20 1580
rect 70 1560 7240 1580
rect 0 1550 7240 1560
rect 5 1545 7240 1550
rect 0 1520 7185 1530
rect 0 1500 20 1520
rect 70 1500 7185 1520
rect 0 1490 7185 1500
rect -305 -6080 -215 1430
rect -85 1235 60 1430
rect -150 135 60 1235
rect 5245 135 5350 1430
rect 6155 135 6260 1430
rect 7145 175 7185 1490
rect -150 -170 -55 135
rect 7145 125 7155 175
rect 7175 125 7185 175
rect 7145 115 7185 125
rect 7200 100 7240 1545
rect 0 90 80 100
rect 0 70 20 90
rect 70 70 80 90
rect 0 60 80 70
rect 7060 60 7240 100
rect 0 30 80 45
rect 0 10 20 30
rect 70 10 80 30
rect 0 0 80 10
rect 7060 40 7185 45
rect 7060 20 7125 40
rect 7175 20 7185 40
rect 7060 5 7185 20
rect 430 -20 7130 -10
rect 430 -40 440 -20
rect 490 -40 1320 -20
rect 1370 -40 2200 -20
rect 2250 -40 3080 -20
rect 3130 -40 3960 -20
rect 4010 -40 4840 -20
rect 4890 -40 5725 -20
rect 5775 -40 6625 -20
rect 6675 -40 7070 -20
rect 7120 -40 7130 -20
rect 430 -50 7130 -40
rect 225 -75 7130 -65
rect 225 -95 235 -75
rect 285 -95 975 -75
rect 1025 -95 1855 -75
rect 1905 -95 2735 -75
rect 2785 -95 3615 -75
rect 3665 -95 4495 -75
rect 4545 -95 5380 -75
rect 5430 -95 6280 -75
rect 6330 -85 7130 -75
rect 6330 -95 7100 -85
rect 225 -105 7100 -95
rect 7090 -135 7100 -105
rect 7120 -135 7130 -85
rect 7090 -145 7130 -135
rect -150 -1465 65 -170
rect 6125 -1465 6230 -170
rect -150 -1770 -55 -1465
rect 0 -1510 85 -1500
rect 0 -1530 20 -1510
rect 70 -1530 85 -1510
rect 0 -1540 85 -1530
rect 7050 -1510 7130 -1500
rect 7050 -1530 7065 -1510
rect 7115 -1530 7130 -1510
rect 7050 -1540 7130 -1530
rect 7145 -1555 7185 5
rect 7200 -1450 7240 60
rect 7280 -20 7350 -10
rect 7280 -40 7290 -20
rect 7340 -40 7350 -20
rect 7280 -50 7350 -40
rect 7200 -1500 7210 -1450
rect 7230 -1500 7240 -1450
rect 7200 -1510 7240 -1500
rect 7255 -115 7295 -105
rect 7255 -165 7265 -115
rect 7285 -165 7295 -115
rect 0 -1570 85 -1555
rect 0 -1590 20 -1570
rect 70 -1590 85 -1570
rect 0 -1600 85 -1590
rect 7060 -1595 7185 -1555
rect 7255 -1535 7295 -165
rect 7255 -1585 7265 -1535
rect 7285 -1585 7295 -1535
rect 7255 -1595 7295 -1585
rect 7310 -1610 7350 -50
rect 430 -1620 7350 -1610
rect 430 -1640 440 -1620
rect 490 -1640 1320 -1620
rect 1370 -1640 2200 -1620
rect 2250 -1640 3080 -1620
rect 3130 -1640 3960 -1620
rect 4010 -1640 4845 -1620
rect 4895 -1640 5725 -1620
rect 5775 -1640 6605 -1620
rect 6655 -1640 7350 -1620
rect 430 -1650 7350 -1640
rect 225 -1675 7295 -1665
rect 225 -1695 235 -1675
rect 285 -1695 975 -1675
rect 1025 -1695 1855 -1675
rect 1905 -1695 2735 -1675
rect 2785 -1695 3615 -1675
rect 3665 -1695 4495 -1675
rect 4545 -1695 5385 -1675
rect 5435 -1695 6245 -1675
rect 6295 -1695 7265 -1675
rect 225 -1705 7265 -1695
rect 7255 -1725 7265 -1705
rect 7285 -1725 7295 -1675
rect -150 -3065 65 -1770
rect -150 -3370 -55 -3065
rect 0 -3110 85 -3100
rect 0 -3130 20 -3110
rect 70 -3130 85 -3110
rect 0 -3140 85 -3130
rect 7255 -3135 7295 -1725
rect 0 -3170 85 -3155
rect 0 -3190 20 -3170
rect 70 -3190 85 -3170
rect 0 -3200 85 -3190
rect 7255 -3185 7265 -3135
rect 7285 -3185 7295 -3135
rect 7255 -3195 7295 -3185
rect 7310 -3210 7350 -1650
rect 430 -3220 7350 -3210
rect 430 -3240 440 -3220
rect 490 -3240 1320 -3220
rect 1370 -3240 2200 -3220
rect 2250 -3240 3080 -3220
rect 3130 -3240 3960 -3220
rect 4010 -3240 4840 -3220
rect 4890 -3240 5720 -3220
rect 5770 -3240 6625 -3220
rect 6675 -3240 7350 -3220
rect 430 -3250 7350 -3240
rect 225 -3275 7295 -3265
rect 225 -3295 235 -3275
rect 285 -3295 975 -3275
rect 1025 -3295 1855 -3275
rect 1905 -3295 2735 -3275
rect 2785 -3295 3615 -3275
rect 3665 -3295 4495 -3275
rect 4545 -3295 5385 -3275
rect 5435 -3295 6260 -3275
rect 6320 -3295 7265 -3275
rect 225 -3305 7265 -3295
rect 7255 -3325 7265 -3305
rect 7285 -3325 7295 -3275
rect -150 -4670 65 -3370
rect 6120 -4670 6240 -3375
rect -150 -4975 -55 -4670
rect 0 -4715 85 -4705
rect 0 -4735 20 -4715
rect 70 -4735 85 -4715
rect 0 -4745 85 -4735
rect 7060 -4740 7220 -4705
rect 7060 -4745 7190 -4740
rect 0 -4775 85 -4760
rect 0 -4795 25 -4775
rect 75 -4795 85 -4775
rect 0 -4805 85 -4795
rect 7060 -4770 7160 -4760
rect 7060 -4790 7100 -4770
rect 7150 -4790 7160 -4770
rect 7060 -4800 7160 -4790
rect 7180 -4790 7190 -4745
rect 7210 -4790 7220 -4740
rect 7180 -4800 7220 -4790
rect 7255 -4740 7295 -3325
rect 7255 -4790 7265 -4740
rect 7285 -4790 7295 -4740
rect 7255 -4800 7295 -4790
rect 7310 -4815 7350 -3250
rect 430 -4825 7350 -4815
rect 430 -4845 440 -4825
rect 490 -4845 1320 -4825
rect 1370 -4845 2200 -4825
rect 2250 -4845 3080 -4825
rect 3130 -4845 3960 -4825
rect 4010 -4845 4840 -4825
rect 4890 -4845 5745 -4825
rect 5795 -4845 6625 -4825
rect 6675 -4845 7350 -4825
rect 430 -4855 7350 -4845
rect 225 -4880 7295 -4870
rect 225 -4900 235 -4880
rect 285 -4900 975 -4880
rect 1025 -4900 1855 -4880
rect 1905 -4900 2735 -4880
rect 2785 -4900 3615 -4880
rect 3665 -4900 4495 -4880
rect 4545 -4900 5400 -4880
rect 5450 -4900 6285 -4880
rect 6330 -4900 7265 -4880
rect 225 -4910 7265 -4900
rect 7120 -4935 7160 -4925
rect -150 -4980 25 -4975
rect -150 -5980 65 -4980
rect -380 -6150 -215 -6080
rect -85 -6140 65 -5980
rect -380 -6385 -315 -6150
rect -150 -6275 65 -6140
rect 5245 -6275 5350 -4980
rect 6150 -6275 6255 -4980
rect 7120 -4985 7130 -4935
rect 7150 -4985 7160 -4935
rect 7120 -6235 7160 -4985
rect -150 -6350 -70 -6275
rect 7120 -6285 7130 -6235
rect 7150 -6285 7160 -6235
rect 7120 -6295 7160 -6285
rect 7180 -4935 7220 -4925
rect 7180 -4985 7190 -4935
rect 7210 -4985 7220 -4935
rect 7180 -6310 7220 -4985
rect 0 -6320 85 -6310
rect 0 -6340 20 -6320
rect 70 -6340 85 -6320
rect 0 -6350 85 -6340
rect 7060 -6345 7220 -6310
rect 7060 -6350 7190 -6345
rect 0 -6380 85 -6365
rect -380 -6475 -260 -6385
rect 0 -6400 20 -6380
rect 70 -6400 85 -6380
rect 0 -6410 85 -6400
rect 7060 -6375 7160 -6365
rect 7060 -6395 7100 -6375
rect 7150 -6395 7160 -6375
rect 7060 -6405 7160 -6395
rect 7180 -6395 7190 -6350
rect 7210 -6395 7220 -6345
rect 7180 -6405 7220 -6395
rect 7255 -4930 7265 -4910
rect 7285 -4930 7295 -4880
rect 7255 -6345 7295 -4930
rect 7255 -6395 7265 -6345
rect 7285 -6395 7295 -6345
rect 7255 -6405 7295 -6395
rect 7310 -6420 7350 -4855
rect 430 -6430 7355 -6420
rect 430 -6450 440 -6430
rect 490 -6450 1320 -6430
rect 1370 -6450 2200 -6430
rect 2250 -6450 3080 -6430
rect 3130 -6450 3960 -6430
rect 4010 -6450 4840 -6430
rect 4890 -6450 5745 -6430
rect 5795 -6450 6625 -6430
rect 6675 -6450 7355 -6430
rect 430 -6460 7355 -6450
rect 225 -6485 7355 -6475
rect 225 -6505 235 -6485
rect 285 -6505 1115 -6485
rect 1165 -6505 1995 -6485
rect 2045 -6505 2875 -6485
rect 2925 -6505 3755 -6485
rect 3805 -6505 4635 -6485
rect 4685 -6505 5540 -6485
rect 5590 -6505 6420 -6485
rect 6470 -6505 7270 -6485
rect 7320 -6505 7355 -6485
rect 225 -6515 7355 -6505
rect 0 -6530 80 -6525
rect 0 -6535 7160 -6530
rect 0 -6555 20 -6535
rect 70 -6540 7160 -6535
rect 70 -6555 7100 -6540
rect 0 -6560 7100 -6555
rect 7150 -6560 7160 -6540
rect 0 -6570 7160 -6560
rect 7180 -6565 7220 -6555
rect 7180 -6585 7190 -6565
rect 0 -6595 7190 -6585
rect 0 -6615 20 -6595
rect 70 -6615 7190 -6595
rect 7210 -6615 7220 -6565
rect 0 -6625 7220 -6615
use dac_unit  dac_unit_0
timestamp 1702614989
transform 1 0 -1115 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_1
timestamp 1702614989
transform 1 0 -235 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_2
timestamp 1702614989
transform 1 0 645 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_3
timestamp 1702614989
transform 1 0 1525 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_4
timestamp 1702614989
transform 1 0 2405 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_5
timestamp 1702614989
transform 1 0 5070 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_6
timestamp 1702614989
transform 1 0 -1115 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_7
timestamp 1702614989
transform 1 0 2405 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_8
timestamp 1702614989
transform 1 0 -235 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_9
timestamp 1702614989
transform 1 0 645 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_10
timestamp 1702614989
transform 1 0 1525 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_11
timestamp 1702614989
transform 1 0 5045 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_12
timestamp 1702614989
transform 1 0 3285 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_13
timestamp 1702614989
transform 1 0 -1115 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_14
timestamp 1702614989
transform 1 0 4165 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_15
timestamp 1702614989
transform 1 0 -235 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_16
timestamp 1702614989
transform 1 0 645 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_17
timestamp 1702614989
transform 1 0 1525 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_18
timestamp 1702614989
transform 1 0 2405 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_19
timestamp 1702614989
transform 1 0 3285 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_20
timestamp 1702614989
transform 1 0 4165 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_21
timestamp 1702614989
transform 1 0 -1115 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_22
timestamp 1702614989
transform 1 0 -235 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_23
timestamp 1702614989
transform 1 0 645 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_24
timestamp 1702614989
transform 1 0 1525 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_25
timestamp 1702614989
transform 1 0 3285 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_26
timestamp 1702614989
transform 1 0 -1115 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_27
timestamp 1702614989
transform 1 0 4165 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_28
timestamp 1702614989
transform 1 0 2405 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_29
timestamp 1702614989
transform 1 0 3285 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_30
timestamp 1702614989
transform 1 0 3285 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_31
timestamp 1702614989
transform 1 0 2405 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_32
timestamp 1702614989
transform 1 0 1525 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_33
timestamp 1702614989
transform 1 0 645 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_34
timestamp 1702614989
transform 1 0 -235 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_35
timestamp 1702614989
transform 1 0 4190 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_36
timestamp 1702614989
transform 1 0 4190 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_37
timestamp 1702614989
transform 1 0 5070 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_38
timestamp 1702614989
transform 1 0 5070 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_40
timestamp 1702614989
transform 1 0 5070 0 1 -50
box 1115 55 2005 1520
use inverter  inverter_0 ~/VLSI_Sine_Gen/layout/dac
timestamp 1693780072
transform 1 0 -40 0 1 -6390
box -240 -145 -30 185
use inverter  inverter_1
timestamp 1693780072
transform 0 1 -220 1 0 1460
box -240 -145 -30 185
use inverter  inverter_2
timestamp 1693780072
transform 0 1 -220 1 0 -140
box -240 -145 -30 185
use inverter  inverter_3
timestamp 1693780072
transform 0 1 -220 1 0 -1740
box -240 -145 -30 185
use inverter  inverter_4
timestamp 1693780072
transform 0 1 -220 1 0 -3340
box -240 -145 -30 185
use inverter  inverter_5
timestamp 1693780072
transform 0 1 -220 1 0 -4945
box -240 -145 -30 185
use inverter  inverter_6
timestamp 1693780072
transform 0 1 -220 1 0 -5910
box -240 -145 -30 185
<< labels >>
rlabel poly 6480 1585 6480 1585 1 Vbp
rlabel poly 6580 1585 6580 1585 1 Vcp
rlabel metal1 7355 -6440 7355 -6440 3 Viout-
rlabel metal1 7355 -6495 7355 -6495 3 Viout+
rlabel metal1 -305 -2540 -305 -2540 7 VN
rlabel metal1 -150 -2280 -150 -2280 7 VP
rlabel locali -415 1570 -415 1570 7 Vphi1
rlabel locali -415 80 -415 80 7 Vphi2
rlabel locali -415 -1520 -415 -1520 7 Vphi3
rlabel locali -415 -3120 -415 -3120 7 Vphi4
rlabel locali -415 -4725 -415 -4725 7 Vphi5
rlabel locali -415 -5880 -415 -5880 7 Vphi6
rlabel locali -380 -6510 -380 -6510 7 Vphi7
<< end >>
