magic
tech sky130A
timestamp 1702365428
<< nmos >>
rect 0 900 50 1500
rect 100 900 150 1500
rect 0 0 50 600
rect 100 0 150 600
<< ndiff >>
rect -50 1485 0 1500
rect -50 915 -35 1485
rect -15 915 0 1485
rect -50 900 0 915
rect 50 1485 100 1500
rect 50 915 65 1485
rect 85 915 100 1485
rect 50 900 100 915
rect 150 1485 200 1500
rect 150 915 165 1485
rect 185 915 200 1485
rect 150 900 200 915
rect -50 585 0 600
rect -50 15 -35 585
rect -15 15 0 585
rect -50 0 0 15
rect 50 585 100 600
rect 50 15 65 585
rect 85 15 100 585
rect 50 0 100 15
rect 150 585 200 600
rect 150 15 165 585
rect 185 15 200 585
rect 150 0 200 15
<< ndiffc >>
rect -35 915 -15 1485
rect 65 915 85 1485
rect 165 915 185 1485
rect -35 15 -15 585
rect 65 15 85 585
rect 165 15 185 585
<< psubdiff >>
rect -100 1490 -50 1500
rect -100 915 -85 1490
rect -65 915 -50 1490
rect -100 900 -50 915
rect -100 590 -50 600
rect -100 15 -85 590
rect -65 15 -50 590
rect -100 0 -50 15
<< psubdiffcont >>
rect -85 915 -65 1490
rect -85 15 -65 590
<< poly >>
rect 0 1500 50 1515
rect 100 1500 150 1515
rect 0 885 50 900
rect 100 885 150 900
rect 0 880 35 885
rect 0 860 5 880
rect 25 860 35 880
rect 0 850 35 860
rect 0 600 50 615
rect 100 600 150 615
rect 0 -15 50 0
rect 100 -15 150 0
rect 0 -20 35 -15
rect 0 -40 5 -20
rect 25 -40 35 -20
rect 0 -50 35 -40
<< polycont >>
rect 5 860 25 880
rect 5 -40 25 -20
<< locali >>
rect -95 1490 -5 1495
rect -95 915 -85 1490
rect -65 1485 -5 1490
rect -65 915 -35 1485
rect -15 915 -5 1485
rect -95 905 -5 915
rect 55 1485 95 1495
rect 55 915 65 1485
rect 85 915 95 1485
rect 55 905 95 915
rect 155 1485 195 1495
rect 155 915 165 1485
rect 185 915 195 1485
rect 155 905 195 915
rect -25 885 -5 905
rect -25 880 35 885
rect -25 865 5 880
rect 0 860 5 865
rect 25 860 35 880
rect 0 850 35 860
rect -95 590 -5 595
rect -95 15 -85 590
rect -65 585 -5 590
rect -65 15 -35 585
rect -15 15 -5 585
rect -95 5 -5 15
rect 55 585 95 595
rect 55 15 65 585
rect 85 15 95 585
rect 55 5 95 15
rect 155 585 195 595
rect 155 15 165 585
rect 185 15 195 585
rect 155 5 195 15
rect -25 -15 -5 5
rect -25 -20 35 -15
rect -25 -35 5 -20
rect 0 -40 5 -35
rect 25 -40 35 -20
rect 0 -50 35 -40
<< end >>
