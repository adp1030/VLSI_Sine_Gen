** sch_path: /home/madvlsi/VLSI_Sine_Gen/simulation/filter/filter_lvs.sch
**.subckt filter_lvs Vout+ Vout- Viout+ Viout-
*.opin Vout+
*.opin Vout-
*.ipin Viout+
*.ipin Viout-
XC3 Vout+ Vout- sky130_fd_pr__cap_mim_m3_1 W=10 L=8 MF=1 m=1
XC4 net1 net2 sky130_fd_pr__cap_mim_m3_1 W=10 L=8 MF=1 m=1
XR7 net2 Vout- GND sky130_fd_pr__res_xhigh_po W=1 L=10 mult=1 m=1
XR8 Viout- net2 GND sky130_fd_pr__res_xhigh_po W=1 L=10 mult=1 m=1
XR9 Vout+ net1 GND sky130_fd_pr__res_xhigh_po W=1 L=10 mult=1 m=1
XR10 net1 Viout+ GND sky130_fd_pr__res_xhigh_po W=1 L=10 mult=1 m=1
XR11 GND Viout- GND sky130_fd_pr__res_xhigh_po W=0.35 L=7 mult=1 m=1
XR12 Viout+ GND GND sky130_fd_pr__res_xhigh_po W=0.35 L=7 mult=1 m=1
**.ends
.GLOBAL GND
.end
