magic
tech sky130A
timestamp 1702370124
<< pdiff >>
rect 295 860 325 960
rect 575 860 605 960
rect 855 860 885 960
rect 1135 860 1165 960
rect 1415 860 1445 960
rect 1695 860 1725 960
rect 1975 860 2005 960
rect 2255 860 2285 960
rect 2535 860 2565 960
rect 2815 860 2845 960
rect 3095 860 3125 960
rect 3375 860 3405 960
rect 3655 860 3685 960
rect 3935 860 3965 960
rect 4215 860 4245 960
rect 295 585 325 685
rect 575 585 605 685
rect 855 585 885 685
rect 1135 585 1165 685
rect 1415 585 1445 685
rect 1695 585 1725 685
rect 1975 585 2005 685
rect 2255 585 2285 685
rect 2535 585 2565 685
rect 2815 585 2845 685
rect 3095 585 3125 685
rect 3375 585 3405 685
rect 3655 585 3685 685
rect 3935 585 3965 685
rect 4215 585 4245 685
<< poly >>
rect -60 895 -20 905
rect -60 875 -50 895
rect -30 875 -20 895
rect -60 865 -20 875
rect 4535 895 4575 905
rect 4535 875 4545 895
rect 4565 875 4575 895
rect 4535 865 4575 875
rect -65 620 -25 630
rect -65 600 -55 620
rect -35 600 -25 620
rect -65 590 -25 600
rect 4540 620 4580 630
rect 4540 600 4550 620
rect 4570 600 4580 620
rect 4540 590 4580 600
<< polycont >>
rect -50 875 -30 895
rect 4545 875 4565 895
rect -55 600 -35 620
rect 4550 600 4570 620
<< locali >>
rect -60 895 -20 905
rect -60 875 -50 895
rect -30 885 -20 895
rect 4535 895 4575 905
rect 4535 885 4545 895
rect -30 875 5 885
rect -60 865 5 875
rect 4510 875 4545 885
rect 4565 875 4575 895
rect 4510 865 4575 875
rect -65 620 -25 630
rect -65 600 -55 620
rect -35 610 -25 620
rect 4540 620 4580 630
rect 4540 610 4550 620
rect -35 600 5 610
rect -65 590 5 600
rect 4510 600 4550 610
rect 4570 600 4580 620
rect 4510 590 4580 600
<< viali >>
rect -50 875 -30 895
rect 4545 875 4565 895
rect -55 600 -35 620
rect 4550 600 4570 620
<< metal1 >>
rect -90 1120 4605 1140
rect -90 625 -70 1120
rect -55 1085 4570 1105
rect -55 895 -25 1085
rect -55 875 -50 895
rect -30 875 -25 895
rect -55 865 -25 875
rect -90 620 -25 625
rect -90 600 -55 620
rect -35 600 -25 620
rect -90 595 -25 600
rect 5 580 25 1050
rect 310 585 330 1055
rect 590 585 610 1055
rect 870 585 890 1055
rect 1150 585 1170 1055
rect 1430 585 1450 1055
rect 1710 585 1730 1055
rect 1990 585 2010 1055
rect 2270 585 2290 1055
rect 2550 585 2570 1055
rect 2830 585 2850 1055
rect 3110 585 3130 1055
rect 3390 585 3410 1055
rect 3670 585 3690 1055
rect 3950 585 3970 1055
rect 4230 585 4250 1055
rect 4540 895 4570 1085
rect 4540 875 4545 895
rect 4565 875 4570 895
rect 4540 865 4570 875
rect 4585 625 4605 1120
rect 4540 620 4605 625
rect 4540 600 4550 620
rect 4570 600 4605 620
rect 4540 595 4605 600
rect 5 70 25 525
rect 310 70 330 530
rect 590 70 610 530
rect 870 70 890 530
rect 1150 70 1170 530
rect 1430 70 1450 530
rect 1710 70 1730 530
rect 1990 70 2010 530
rect 2270 70 2290 530
rect 2550 70 2570 530
rect 2830 70 2850 530
rect 3110 70 3130 530
rect 3390 70 3410 530
rect 3670 70 3690 530
rect 3950 70 3970 530
rect 4230 70 4250 530
rect 5 0 25 40
rect 310 0 330 40
rect 590 0 610 40
rect 870 0 890 40
rect 1150 0 1170 40
rect 1430 0 1450 40
rect 1710 0 1730 40
rect 1990 0 2010 40
rect 2270 0 2290 40
rect 2550 0 2570 40
rect 2830 0 2850 40
rect 3110 0 3130 40
rect 3390 0 3410 40
rect 3670 0 3690 40
rect 3950 0 3970 40
rect 4230 0 4250 40
use csrl_dff1  csrl_dff1_0 ~/VLSI_Sine_Gen/layout/shift_register
timestamp 1702367094
transform 1 0 550 0 1 270
box -565 -270 -220 805
use csrl_dff2  csrl_dff2_0 ~/VLSI_Sine_Gen/layout/shift_register
timestamp 1702366369
transform 1 0 830 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_1
timestamp 1702366369
transform 1 0 1110 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_2
timestamp 1702366369
transform 1 0 1390 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_3
timestamp 1702366369
transform 1 0 1670 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_4
timestamp 1702366369
transform 1 0 1950 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_5
timestamp 1702366369
transform 1 0 2230 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_6
timestamp 1702366369
transform 1 0 2510 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_7
timestamp 1702366369
transform 1 0 2790 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_8
timestamp 1702366369
transform 1 0 3070 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_9
timestamp 1702366369
transform 1 0 3350 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_10
timestamp 1702366369
transform 1 0 3630 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_11
timestamp 1702366369
transform 1 0 3910 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_12
timestamp 1702366369
transform 1 0 4190 0 1 270
box -540 -270 -220 805
use csrl_dff2  csrl_dff2_13
timestamp 1702366369
transform 1 0 4470 0 1 270
box -540 -270 -220 805
use csrl_dff3  csrl_dff3_0 ~/VLSI_Sine_Gen/layout/shift_register
timestamp 1702367186
transform 1 0 4750 0 1 270
box -540 -270 -220 805
<< end >>
