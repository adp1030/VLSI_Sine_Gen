magic
tech sky130A
timestamp 1702709769
<< psubdiff >>
rect 1450 3200 1600 3215
rect 1450 3170 1465 3200
rect 1585 3170 1600 3200
rect 1450 3155 1600 3170
rect 730 1830 880 1845
rect 730 1800 745 1830
rect 865 1800 880 1830
rect 730 1785 880 1800
rect 630 1035 690 1050
rect 630 915 645 1035
rect 675 915 690 1035
rect 630 900 690 915
rect 1450 630 1510 645
rect 1450 510 1465 630
rect 1495 510 1510 630
rect 1450 495 1510 510
<< psubdiffcont >>
rect 1465 3170 1585 3200
rect 745 1800 865 1830
rect 645 915 675 1035
rect 1465 510 1495 630
<< xpolycontact >>
rect 610 3190 830 3225
rect 1180 3190 1400 3225
rect 610 3130 830 3165
rect 1180 3130 1400 3165
rect 730 3015 950 3050
rect 1300 3015 1520 3050
rect 730 2910 950 2945
rect 1300 2910 1520 2945
rect 715 1700 935 1735
rect 1285 1700 1505 1735
rect 545 1225 580 1445
rect 545 655 580 875
rect 610 610 830 645
rect 1180 610 1400 645
rect 610 550 830 585
rect 1180 550 1400 585
<< xpolyres >>
rect 830 3190 1180 3225
rect 830 3130 1180 3165
rect 950 3015 1300 3050
rect 950 2910 1300 2945
rect 935 1700 1285 1735
rect 545 875 580 1225
rect 830 610 1180 645
rect 830 550 1180 585
<< locali >>
rect 680 3270 830 3285
rect 680 3240 695 3270
rect 815 3240 830 3270
rect 680 3225 830 3240
rect 1180 3165 1400 3190
rect 1455 3200 1595 3210
rect 1455 3170 1465 3200
rect 1585 3170 1595 3200
rect 1455 3160 1595 3170
rect 610 3110 830 3130
rect 535 3085 1520 3110
rect 1300 3050 1520 3085
rect 730 3000 950 3015
rect 730 2990 880 3000
rect 730 2960 745 2990
rect 865 2960 880 2990
rect 730 2945 880 2960
rect 1520 2910 1685 2945
rect 1595 2840 1675 2910
rect 1595 2740 1610 2840
rect 1660 2740 1675 2840
rect 1595 2725 1675 2740
rect 1595 2045 1675 2060
rect 1595 1945 1610 2045
rect 1660 1945 1675 2045
rect 735 1830 875 1840
rect 735 1800 745 1830
rect 865 1800 875 1830
rect 735 1790 875 1800
rect 1595 1735 1675 1945
rect 545 1700 715 1735
rect 1505 1700 1685 1735
rect 545 1655 580 1700
rect 545 1640 625 1655
rect 545 1540 560 1640
rect 610 1540 625 1640
rect 545 1525 625 1540
rect 1600 1640 1680 1655
rect 1600 1540 1615 1640
rect 1665 1540 1680 1640
rect 1600 1525 1680 1540
rect 545 1445 580 1525
rect 635 1035 685 1045
rect 635 915 645 1035
rect 675 915 685 1035
rect 635 905 685 915
rect 545 645 580 655
rect 535 610 610 645
rect 1180 585 1400 610
rect 1455 630 1505 640
rect 680 535 830 550
rect 680 505 695 535
rect 815 505 830 535
rect 680 490 830 505
rect 1455 510 1465 630
rect 1495 510 1505 630
rect 1455 500 1505 510
<< viali >>
rect 695 3240 815 3270
rect 1465 3170 1585 3200
rect 745 2960 865 2990
rect 1610 2740 1660 2840
rect 1610 1945 1660 2045
rect 745 1800 865 1830
rect 560 1540 610 1640
rect 1615 1540 1665 1640
rect 645 915 675 1035
rect 695 505 815 535
rect 1465 510 1495 630
<< metal1 >>
rect 650 3270 1630 3285
rect 650 3240 695 3270
rect 815 3240 1630 3270
rect 650 3200 1630 3240
rect 650 3170 1465 3200
rect 1585 3170 1630 3200
rect 650 3100 1630 3170
rect 650 1855 690 3100
rect 730 2990 880 3005
rect 730 2960 745 2990
rect 865 2960 880 2990
rect 730 2945 880 2960
rect 1595 2840 1675 2855
rect 1595 2740 1610 2840
rect 1660 2740 1675 2840
rect 1595 2725 1675 2740
rect 1595 2045 1675 2060
rect 1595 1945 1610 2045
rect 1660 1945 1675 2045
rect 1595 1930 1675 1945
rect 650 1830 915 1855
rect 650 1800 745 1830
rect 865 1800 915 1830
rect 650 1765 915 1800
rect 545 1640 625 1655
rect 545 1540 560 1640
rect 610 1540 625 1640
rect 545 1525 625 1540
rect 650 1475 690 1765
rect 1600 1640 1680 1655
rect 1600 1540 1615 1640
rect 1665 1540 1680 1640
rect 1600 1525 1680 1540
rect 630 1035 690 1475
rect 630 915 645 1035
rect 675 915 690 1035
rect 630 650 690 915
rect 630 630 1525 650
rect 630 550 1465 630
rect 535 535 1465 550
rect 535 505 695 535
rect 815 510 1465 535
rect 1495 510 1525 630
rect 815 505 1525 510
rect 535 490 1525 505
<< via1 >>
rect 745 2960 865 2990
rect 1610 2740 1660 2840
rect 1610 1945 1660 2045
rect 560 1540 610 1640
rect 1615 1540 1665 1640
<< metal2 >>
rect 730 2990 880 3005
rect 730 2960 745 2990
rect 865 2975 880 2990
rect 865 2960 1575 2975
rect 730 2945 1575 2960
rect 1545 1655 1575 2945
rect 1595 2840 1675 2855
rect 1595 2740 1610 2840
rect 1660 2740 1675 2840
rect 1595 2725 1675 2740
rect 1595 2045 1675 2060
rect 1595 1945 1610 2045
rect 1660 1945 1675 2045
rect 1595 1930 1675 1945
rect 545 1640 625 1655
rect 545 1540 560 1640
rect 610 1540 625 1640
rect 545 1525 625 1540
rect 1545 1640 1680 1655
rect 1545 1540 1615 1640
rect 1665 1540 1680 1640
rect 1545 1525 1680 1540
<< via2 >>
rect 1610 2740 1660 2840
rect 1610 1945 1660 2045
rect 560 1540 610 1640
rect 1615 1540 1665 1640
<< metal3 >>
rect 690 2060 1530 2890
rect 1595 2840 1675 2855
rect 1595 2740 1610 2840
rect 1660 2740 1675 2840
rect 1595 2725 1675 2740
rect 690 2045 1675 2060
rect 690 1945 1610 2045
rect 1660 1945 1675 2045
rect 690 1930 1675 1945
rect 690 1850 1530 1930
rect 700 1655 1530 1685
rect 545 1640 1530 1655
rect 545 1540 560 1640
rect 610 1540 1530 1640
rect 545 1525 1530 1540
rect 1600 1640 1680 1655
rect 1600 1540 1615 1640
rect 1665 1540 1680 1640
rect 1600 1525 1680 1540
rect 700 655 1530 1525
<< via3 >>
rect 1610 2740 1660 2840
rect 1615 1540 1665 1640
<< mimcap >>
rect 710 2840 1510 2870
rect 710 2740 1400 2840
rect 1480 2740 1510 2840
rect 710 1870 1510 2740
rect 715 1640 1515 1670
rect 715 1540 1405 1640
rect 1485 1540 1515 1640
rect 715 670 1515 1540
<< mimcapcontact >>
rect 1400 2740 1480 2840
rect 1405 1540 1485 1640
<< metal4 >>
rect 1385 2840 1675 2855
rect 1385 2740 1400 2840
rect 1480 2740 1610 2840
rect 1660 2740 1675 2840
rect 1385 2725 1675 2740
rect 1390 1640 1680 1655
rect 1390 1540 1405 1640
rect 1485 1540 1615 1640
rect 1665 1540 1680 1640
rect 1390 1525 1680 1540
<< labels >>
rlabel locali 1685 2930 1685 2930 3 Vout+
rlabel locali 1685 1720 1685 1720 3 Vout-
rlabel locali 535 625 535 625 7 Viout-
rlabel metal1 535 520 535 520 7 VN
rlabel locali 535 3100 535 3100 7 Viout+
<< end >>
