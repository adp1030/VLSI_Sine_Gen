magic
tech sky130A
timestamp 1702614989
<< nwell >>
rect 1115 155 2005 1510
<< pmos >>
rect 1185 885 1235 1485
rect 1385 885 1435 1485
rect 1485 885 1535 1485
rect 1585 885 1635 1485
rect 1685 885 1735 1485
rect 1885 885 1935 1485
rect 1285 180 1335 780
rect 1385 180 1435 780
rect 1485 180 1535 780
rect 1585 180 1635 780
rect 1685 180 1735 780
rect 1785 180 1835 780
<< pdiff >>
rect 1135 1470 1185 1485
rect 1135 900 1150 1470
rect 1170 900 1185 1470
rect 1135 885 1185 900
rect 1235 1470 1285 1485
rect 1335 1470 1385 1485
rect 1235 900 1250 1470
rect 1270 900 1285 1470
rect 1335 900 1350 1470
rect 1370 900 1385 1470
rect 1235 885 1285 900
rect 1335 885 1385 900
rect 1435 1470 1485 1485
rect 1435 900 1450 1470
rect 1470 900 1485 1470
rect 1435 885 1485 900
rect 1535 1470 1585 1485
rect 1535 900 1550 1470
rect 1570 900 1585 1470
rect 1535 885 1585 900
rect 1635 1470 1685 1485
rect 1635 900 1650 1470
rect 1670 900 1685 1470
rect 1635 885 1685 900
rect 1735 1470 1785 1485
rect 1835 1470 1885 1485
rect 1735 900 1750 1470
rect 1770 900 1785 1470
rect 1835 900 1850 1470
rect 1870 900 1885 1470
rect 1735 885 1785 900
rect 1835 885 1885 900
rect 1935 1470 1985 1485
rect 1935 900 1950 1470
rect 1970 900 1985 1470
rect 1935 885 1985 900
rect 1235 765 1285 780
rect 1235 195 1250 765
rect 1270 195 1285 765
rect 1235 180 1285 195
rect 1335 765 1385 780
rect 1335 195 1350 765
rect 1370 195 1385 765
rect 1335 180 1385 195
rect 1435 765 1485 780
rect 1435 195 1450 765
rect 1470 195 1485 765
rect 1435 180 1485 195
rect 1535 765 1585 780
rect 1535 195 1550 765
rect 1570 195 1585 765
rect 1535 180 1585 195
rect 1635 765 1685 780
rect 1635 195 1650 765
rect 1670 195 1685 765
rect 1635 180 1685 195
rect 1735 765 1785 780
rect 1735 195 1750 765
rect 1770 195 1785 765
rect 1735 180 1785 195
rect 1835 765 1885 780
rect 1835 195 1850 765
rect 1870 195 1885 765
rect 1835 180 1885 195
<< pdiffc >>
rect 1150 900 1170 1470
rect 1250 900 1270 1470
rect 1350 900 1370 1470
rect 1450 900 1470 1470
rect 1550 900 1570 1470
rect 1650 900 1670 1470
rect 1750 900 1770 1470
rect 1850 900 1870 1470
rect 1950 900 1970 1470
rect 1250 195 1270 765
rect 1350 195 1370 765
rect 1450 195 1470 765
rect 1550 195 1570 765
rect 1650 195 1670 765
rect 1750 195 1770 765
rect 1850 195 1870 765
<< nsubdiff >>
rect 1285 1470 1335 1485
rect 1285 900 1300 1470
rect 1320 900 1335 1470
rect 1285 885 1335 900
rect 1785 1470 1835 1485
rect 1785 900 1800 1470
rect 1820 900 1835 1470
rect 1785 885 1835 900
rect 1185 765 1235 780
rect 1185 195 1200 765
rect 1220 195 1235 765
rect 1185 180 1235 195
rect 1885 765 1935 780
rect 1885 195 1900 765
rect 1920 195 1935 765
rect 1885 180 1935 195
<< nsubdiffcont >>
rect 1300 900 1320 1470
rect 1800 900 1820 1470
rect 1200 195 1220 765
rect 1900 195 1920 765
<< poly >>
rect 1185 1485 1235 1505
rect 1385 1485 1435 1520
rect 1485 1505 1635 1520
rect 1485 1485 1535 1505
rect 1585 1485 1635 1505
rect 1685 1485 1735 1505
rect 1885 1485 1935 1505
rect 1185 865 1235 885
rect 1185 855 1280 865
rect 1185 850 1250 855
rect 1240 835 1250 850
rect 1270 835 1280 855
rect 1240 825 1280 835
rect 1385 840 1435 885
rect 1485 865 1535 885
rect 1585 865 1635 885
rect 1685 840 1735 885
rect 1885 865 1935 885
rect 1385 825 1735 840
rect 1840 855 1935 865
rect 1840 835 1850 855
rect 1870 850 1935 855
rect 1870 835 1880 850
rect 1840 825 1880 835
rect 1285 780 1335 800
rect 1385 780 1435 800
rect 1485 780 1535 800
rect 1585 780 1635 800
rect 1685 780 1735 800
rect 1785 780 1835 800
rect 1285 165 1335 180
rect 1240 155 1335 165
rect 1240 135 1250 155
rect 1270 150 1335 155
rect 1270 135 1280 150
rect 1240 125 1280 135
rect 1385 85 1435 180
rect 1485 140 1535 180
rect 1485 120 1495 140
rect 1515 120 1535 140
rect 1485 110 1535 120
rect 1585 140 1635 180
rect 1585 120 1605 140
rect 1625 120 1635 140
rect 1585 110 1635 120
rect 1385 65 1405 85
rect 1425 65 1435 85
rect 1385 55 1435 65
rect 1685 85 1735 180
rect 1785 165 1835 180
rect 1785 155 1880 165
rect 1785 150 1850 155
rect 1840 135 1850 150
rect 1870 135 1880 155
rect 1840 125 1880 135
rect 1685 65 1695 85
rect 1715 65 1735 85
rect 1685 55 1735 65
<< polycont >>
rect 1250 835 1270 855
rect 1850 835 1870 855
rect 1250 135 1270 155
rect 1495 120 1515 140
rect 1605 120 1625 140
rect 1405 65 1425 85
rect 1850 135 1870 155
rect 1695 65 1715 85
<< locali >>
rect 1140 1500 1480 1520
rect 1140 1470 1180 1500
rect 1140 900 1150 1470
rect 1170 900 1180 1470
rect 1140 890 1180 900
rect 1240 1470 1380 1480
rect 1240 900 1250 1470
rect 1270 900 1300 1470
rect 1320 900 1350 1470
rect 1370 900 1380 1470
rect 1240 890 1380 900
rect 1440 1470 1480 1500
rect 1640 1500 1980 1520
rect 1440 900 1450 1470
rect 1470 900 1480 1470
rect 1440 890 1480 900
rect 1540 1470 1580 1480
rect 1540 900 1550 1470
rect 1570 900 1580 1470
rect 1240 855 1280 890
rect 1240 835 1250 855
rect 1270 835 1280 855
rect 1240 825 1280 835
rect 1340 840 1420 850
rect 1340 820 1350 840
rect 1410 820 1420 840
rect 1540 830 1580 900
rect 1640 1470 1680 1500
rect 1640 900 1650 1470
rect 1670 900 1680 1470
rect 1640 890 1680 900
rect 1740 1470 1880 1480
rect 1740 900 1750 1470
rect 1770 900 1800 1470
rect 1820 900 1850 1470
rect 1870 900 1880 1470
rect 1740 890 1880 900
rect 1940 1470 1980 1500
rect 1940 900 1950 1470
rect 1970 900 1980 1470
rect 1940 890 1980 900
rect 1840 855 1880 890
rect 1700 840 1780 850
rect 1340 810 1420 820
rect 1190 765 1280 775
rect 1190 195 1200 765
rect 1220 195 1250 765
rect 1270 195 1280 765
rect 1190 185 1280 195
rect 1240 155 1280 185
rect 1240 135 1250 155
rect 1270 135 1280 155
rect 1240 125 1280 135
rect 1340 765 1380 810
rect 1340 195 1350 765
rect 1370 195 1380 765
rect 1340 185 1380 195
rect 1440 795 1680 830
rect 1700 820 1710 840
rect 1770 820 1780 840
rect 1840 835 1850 855
rect 1870 835 1880 855
rect 1840 825 1880 835
rect 1700 810 1780 820
rect 1440 765 1480 795
rect 1440 195 1450 765
rect 1470 195 1480 765
rect 1440 185 1480 195
rect 1540 765 1580 775
rect 1540 195 1550 765
rect 1570 195 1580 765
rect 1540 185 1580 195
rect 1640 765 1680 795
rect 1640 195 1650 765
rect 1670 195 1680 765
rect 1640 185 1680 195
rect 1740 765 1780 810
rect 1740 195 1750 765
rect 1770 195 1780 765
rect 1740 185 1780 195
rect 1840 765 1930 775
rect 1840 195 1850 765
rect 1870 195 1900 765
rect 1920 195 1930 765
rect 1840 185 1930 195
rect 1340 55 1375 185
rect 1485 140 1525 150
rect 1485 120 1495 140
rect 1515 120 1525 140
rect 1485 110 1525 120
rect 1395 85 1435 95
rect 1395 65 1405 85
rect 1425 65 1435 85
rect 1395 55 1435 65
rect 1545 55 1575 185
rect 1840 155 1880 185
rect 1595 140 1635 150
rect 1595 120 1605 140
rect 1625 120 1635 140
rect 1840 135 1850 155
rect 1870 135 1880 155
rect 1840 125 1880 135
rect 1595 110 1635 120
rect 1685 85 1725 95
rect 1685 65 1695 85
rect 1715 65 1725 85
rect 1685 55 1725 65
<< viali >>
rect 1250 900 1270 1470
rect 1300 900 1320 1470
rect 1350 900 1370 1470
rect 1350 820 1410 840
rect 1750 900 1770 1470
rect 1800 900 1820 1470
rect 1850 900 1870 1470
rect 1200 195 1220 765
rect 1250 195 1270 765
rect 1710 820 1770 840
rect 1850 195 1870 765
rect 1900 195 1920 765
rect 1495 120 1515 140
rect 1405 65 1425 85
rect 1605 120 1625 140
rect 1695 65 1715 85
<< metal1 >>
rect 1135 1480 1985 1485
rect 1115 1470 2005 1480
rect 1115 900 1250 1470
rect 1270 900 1300 1470
rect 1320 900 1350 1470
rect 1370 900 1750 1470
rect 1770 900 1800 1470
rect 1820 900 1850 1470
rect 1870 900 2005 1470
rect 1115 885 2005 900
rect 1115 780 1305 885
rect 1340 840 1780 850
rect 1340 820 1350 840
rect 1410 820 1710 840
rect 1770 820 1780 840
rect 1340 810 1780 820
rect 1815 780 2005 885
rect 1115 765 2005 780
rect 1115 195 1200 765
rect 1220 195 1250 765
rect 1270 195 1850 765
rect 1870 195 1900 765
rect 1920 195 2005 765
rect 1115 185 2005 195
rect 1185 180 1935 185
rect 1115 140 2005 150
rect 1115 120 1495 140
rect 1515 120 1605 140
rect 1625 120 2005 140
rect 1115 110 2005 120
rect 1115 85 2005 95
rect 1115 65 1405 85
rect 1425 65 1695 85
rect 1715 65 2005 85
rect 1115 55 2005 65
<< labels >>
rlabel poly 1510 1520 1510 1520 1 Vcp
port 2 n
rlabel poly 1410 1520 1410 1520 1 Vbp
port 1 n
rlabel metal1 1115 1180 1115 1180 7 VP
port 7 w
rlabel metal1 1115 130 1115 130 7 Vphi
port 3 w
rlabel metal1 1115 75 1115 75 7 Vphi_b
port 4 w
rlabel locali 1560 55 1560 55 5 Viun
port 6 s
rlabel locali 1360 55 1360 55 5 Viup
port 5 s
<< end >>
