magic
tech sky130A
timestamp 1695756208
<< nwell >>
rect -50 295 290 810
<< nmos >>
rect 10 -140 25 260
rect 75 160 90 260
rect 140 160 155 260
rect 205 160 220 260
rect 75 -105 90 -5
rect 140 -105 155 -5
rect 205 -105 220 -5
<< pmos >>
rect 20 615 35 715
rect 85 615 100 715
rect 20 315 35 415
rect 85 315 100 415
rect 150 315 165 715
rect 205 560 220 660
rect 205 315 220 415
<< ndiff >>
rect -40 240 10 260
rect -40 180 -25 240
rect -5 180 10 240
rect -40 160 10 180
rect -20 -40 10 160
rect -40 -60 10 -40
rect -40 -120 -25 -60
rect -5 -120 10 -60
rect -40 -140 10 -120
rect 25 160 75 260
rect 90 245 140 260
rect 90 175 105 245
rect 125 175 140 245
rect 90 160 140 175
rect 155 245 205 260
rect 155 175 170 245
rect 190 175 205 245
rect 155 160 205 175
rect 220 245 270 260
rect 220 175 235 245
rect 255 175 270 245
rect 220 160 270 175
rect 25 -5 55 160
rect 25 -105 75 -5
rect 90 -20 140 -5
rect 90 -90 105 -20
rect 125 -90 140 -20
rect 90 -105 140 -90
rect 155 -20 205 -5
rect 155 -90 170 -20
rect 190 -90 205 -20
rect 155 -105 205 -90
rect 220 -20 270 -5
rect 220 -90 235 -20
rect 255 -90 270 -20
rect 220 -105 270 -90
rect 25 -140 55 -105
<< pdiff >>
rect -30 700 20 715
rect -30 630 -15 700
rect 5 630 20 700
rect -30 615 20 630
rect 35 700 85 715
rect 35 630 50 700
rect 70 630 85 700
rect 35 615 85 630
rect 100 700 150 715
rect 100 630 115 700
rect 135 630 150 700
rect 100 615 150 630
rect 125 415 150 615
rect -30 400 20 415
rect -30 330 -15 400
rect 5 330 20 400
rect -30 315 20 330
rect 35 400 85 415
rect 35 330 50 400
rect 70 330 85 400
rect 35 315 85 330
rect 100 400 150 415
rect 100 330 115 400
rect 135 330 150 400
rect 100 315 150 330
rect 165 660 190 715
rect 165 560 205 660
rect 220 645 270 660
rect 220 575 235 645
rect 255 575 270 645
rect 220 560 270 575
rect 165 415 190 560
rect 165 315 205 415
rect 220 400 270 415
rect 220 330 235 400
rect 255 330 270 400
rect 220 315 270 330
<< ndiffc >>
rect -25 180 -5 240
rect -25 -120 -5 -60
rect 105 175 125 245
rect 170 175 190 245
rect 235 175 255 245
rect 105 -90 125 -20
rect 170 -90 190 -20
rect 235 -90 255 -20
<< pdiffc >>
rect -15 630 5 700
rect 50 630 70 700
rect 115 630 135 700
rect -15 330 5 400
rect 50 330 70 400
rect 115 330 135 400
rect 235 575 255 645
rect 235 330 255 400
<< psubdiff >>
rect 155 -155 270 -140
rect 155 -175 175 -155
rect 250 -175 270 -155
rect 155 -190 270 -175
<< nsubdiff >>
rect 220 770 270 790
rect 220 705 235 770
rect 255 705 270 770
rect 220 690 270 705
<< psubdiffcont >>
rect 175 -175 250 -155
<< nsubdiffcont >>
rect 235 705 255 770
<< poly >>
rect 20 715 35 730
rect 85 715 100 730
rect 150 715 165 730
rect 20 605 35 615
rect -35 590 35 605
rect -35 440 -20 590
rect 85 560 100 615
rect 5 550 45 560
rect 5 530 15 550
rect 35 530 45 550
rect 5 520 45 530
rect 70 550 110 560
rect 70 530 80 550
rect 100 530 110 550
rect 70 520 110 530
rect 25 480 40 520
rect 25 465 100 480
rect -35 425 35 440
rect 20 415 35 425
rect 85 415 100 465
rect 205 660 220 675
rect 205 545 220 560
rect 205 535 245 545
rect 205 515 215 535
rect 235 515 245 535
rect 205 505 245 515
rect 225 465 265 475
rect 225 450 235 465
rect 205 445 235 450
rect 255 445 265 465
rect 205 435 265 445
rect 205 415 220 435
rect 20 300 35 315
rect 85 300 100 315
rect 150 300 165 315
rect 10 285 35 300
rect 75 285 100 300
rect 140 285 165 300
rect 10 260 25 285
rect 75 260 90 285
rect 140 260 155 285
rect 205 260 220 315
rect 75 145 90 160
rect 75 135 115 145
rect 75 115 85 135
rect 105 115 115 135
rect 75 105 115 115
rect 65 70 105 80
rect 65 50 75 70
rect 95 50 105 70
rect 65 40 105 50
rect 75 -5 90 40
rect 140 -5 155 160
rect 205 145 220 160
rect 205 135 285 145
rect 205 130 255 135
rect 245 115 255 130
rect 275 115 285 135
rect 245 105 285 115
rect 180 95 220 105
rect 180 75 190 95
rect 210 75 220 95
rect 180 65 220 75
rect 205 -5 220 65
rect 75 -120 90 -105
rect 140 -115 155 -105
rect 130 -130 155 -115
rect 205 -120 220 -105
rect 10 -220 25 -140
rect 130 -220 145 -130
rect 10 -230 50 -220
rect 10 -250 20 -230
rect 40 -250 50 -230
rect 10 -260 50 -250
rect 130 -230 170 -220
rect 130 -250 140 -230
rect 160 -250 170 -230
rect 130 -260 170 -250
<< polycont >>
rect 15 530 35 550
rect 80 530 100 550
rect 215 515 235 535
rect 235 445 255 465
rect 85 115 105 135
rect 75 50 95 70
rect 255 115 275 135
rect 190 75 210 95
rect 20 -250 40 -230
rect 140 -250 160 -230
<< locali >>
rect 225 770 265 785
rect 225 750 235 770
rect 125 730 235 750
rect 125 710 145 730
rect -25 700 15 710
rect -25 640 -15 700
rect -50 630 -15 640
rect 5 630 15 700
rect -50 620 15 630
rect 40 700 80 710
rect 40 630 50 700
rect 70 630 80 700
rect 40 620 80 630
rect 105 700 145 710
rect 105 630 115 700
rect 135 630 145 700
rect 225 705 235 730
rect 255 705 265 770
rect 225 695 265 705
rect 105 620 145 630
rect 225 645 265 655
rect 40 600 60 620
rect 25 580 60 600
rect 25 560 45 580
rect 225 575 235 645
rect 255 640 265 645
rect 255 620 290 640
rect 255 585 265 620
rect 255 575 285 585
rect 225 565 285 575
rect 5 550 45 560
rect 5 530 15 550
rect 35 530 45 550
rect 5 520 45 530
rect 70 550 110 560
rect 70 530 80 550
rect 100 530 110 550
rect 205 535 245 545
rect 205 530 215 535
rect 70 520 110 530
rect 70 500 90 520
rect 60 480 90 500
rect 180 515 215 530
rect 235 515 245 535
rect 180 505 245 515
rect 60 410 80 480
rect 180 410 200 505
rect 265 475 285 565
rect 225 465 285 475
rect 225 445 235 465
rect 255 455 285 465
rect 255 445 265 455
rect 225 435 265 445
rect -25 400 15 410
rect -25 340 -15 400
rect -50 330 -15 340
rect 5 330 15 400
rect -50 320 15 330
rect 40 400 80 410
rect 40 330 50 400
rect 70 330 80 400
rect 40 320 80 330
rect 105 400 145 410
rect 105 330 115 400
rect 135 330 145 400
rect 105 320 145 330
rect 180 400 265 410
rect 180 390 235 400
rect 60 255 80 320
rect 180 255 200 390
rect 225 330 235 390
rect 255 340 265 400
rect 255 330 290 340
rect 225 320 290 330
rect -35 240 5 255
rect -35 180 -25 240
rect -5 180 5 240
rect -35 165 5 180
rect 35 245 135 255
rect 35 235 105 245
rect 35 80 55 235
rect 95 175 105 235
rect 125 175 135 245
rect 95 165 135 175
rect 160 245 200 255
rect 160 175 170 245
rect 190 175 200 245
rect 160 165 200 175
rect 225 245 265 255
rect 225 175 235 245
rect 255 175 265 245
rect 225 165 265 175
rect 75 135 115 145
rect 75 115 85 135
rect 105 125 115 135
rect 105 115 150 125
rect 75 105 150 115
rect 35 70 105 80
rect 35 60 75 70
rect 65 50 75 60
rect 95 50 105 70
rect 65 40 105 50
rect 130 25 150 105
rect 180 105 200 165
rect 245 135 285 145
rect 245 115 255 135
rect 275 115 285 135
rect 245 105 285 115
rect 180 95 220 105
rect 180 75 190 95
rect 210 75 220 95
rect 180 65 220 75
rect 245 45 265 105
rect 115 5 150 25
rect 180 25 265 45
rect 115 -10 135 5
rect 180 -10 200 25
rect 95 -20 135 -10
rect -35 -60 5 -45
rect -35 -120 -25 -60
rect -5 -120 5 -60
rect 95 -90 105 -20
rect 125 -90 135 -20
rect 95 -100 135 -90
rect 160 -20 200 -10
rect 160 -90 170 -20
rect 190 -90 200 -20
rect 160 -100 200 -90
rect 225 -20 265 -10
rect 225 -90 235 -20
rect 255 -90 265 -20
rect 225 -100 265 -90
rect -35 -135 5 -120
rect 225 -145 245 -100
rect 160 -155 265 -145
rect 160 -175 175 -155
rect 250 -175 265 -155
rect 160 -185 265 -175
rect 10 -230 50 -220
rect 10 -250 20 -230
rect 40 -250 50 -230
rect 10 -260 50 -250
rect 130 -230 170 -220
rect 130 -250 140 -230
rect 160 -250 170 -230
rect 130 -260 170 -250
<< viali >>
rect 115 630 135 700
rect 235 705 255 770
rect 115 330 135 400
rect -25 180 -5 240
rect 235 175 255 245
rect -25 -120 -5 -60
rect 235 -90 255 -20
rect 175 -175 250 -155
rect 20 -250 40 -230
rect 140 -250 160 -230
<< metal1 >>
rect -50 770 290 790
rect -50 705 235 770
rect 255 705 290 770
rect -50 700 290 705
rect -50 630 115 700
rect 135 630 290 700
rect -50 400 290 630
rect -50 330 115 400
rect 135 330 290 400
rect -50 315 290 330
rect -50 245 290 260
rect -50 240 235 245
rect -50 180 -25 240
rect -5 180 235 240
rect -50 175 235 180
rect 255 175 290 245
rect -50 -20 290 175
rect -50 -60 235 -20
rect -50 -120 -25 -60
rect -5 -90 235 -60
rect 255 -90 290 -20
rect -5 -120 290 -90
rect -50 -155 290 -120
rect -50 -175 175 -155
rect 250 -175 290 -155
rect -50 -190 290 -175
rect -50 -230 290 -220
rect -50 -250 20 -230
rect 40 -250 140 -230
rect 160 -250 290 -230
rect -50 -260 290 -250
<< labels >>
rlabel metal1 -50 50 -50 50 3 VN
port 7 e
rlabel locali -50 330 -50 330 7 DB
port 2 w
rlabel metal1 -50 -240 -50 -240 7 CLK
port 3 w
rlabel metal1 -50 560 -50 560 7 VP
port 6 w
rlabel locali -50 630 -50 630 7 D
port 1 w
rlabel locali 290 330 290 330 3 QB
port 5 e
rlabel locali 290 630 290 630 3 Q
port 4 e
<< end >>
