magic
tech sky130A
timestamp 1702887642
<< poly >>
rect -4525 8810 -4510 8820
rect -4980 8795 -4510 8810
rect -4815 8090 -4775 8100
rect -4815 8075 -4805 8090
rect -5010 8070 -4805 8075
rect -4785 8070 -4775 8090
rect -5010 8060 -4775 8070
<< polycont >>
rect -4805 8070 -4785 8090
<< locali >>
rect -4530 8735 -4090 8775
rect -4885 7385 -4865 8485
rect -4815 8090 -4775 8100
rect -4815 8070 -4805 8090
rect -4785 8080 -4775 8090
rect -4530 8080 -4510 8735
rect -4785 8070 -4510 8080
rect -4815 8060 -4510 8070
rect -7290 7365 -7060 7385
rect -5000 7365 -4865 7385
rect -5990 7080 -5950 7090
rect -5990 7030 -5980 7080
rect -5960 7030 -5950 7080
rect -5990 6935 -5950 7030
rect -5990 6925 -5910 6935
rect -5990 6905 -5980 6925
rect -5920 6905 -5910 6925
rect -5990 6895 -5910 6905
rect -5000 6620 -4980 7365
rect -5660 6600 -5425 6620
rect -5075 6600 -4980 6620
rect -4960 6865 -4915 6905
rect -5660 6325 -5465 6345
rect -5485 6250 -5465 6325
rect -4960 6270 -4940 6865
rect -5070 6250 -4940 6270
rect -5660 6050 -5510 6070
rect -5530 5920 -5510 6050
rect -5530 5900 -5425 5920
rect -5075 5900 -4905 5920
rect -5660 5775 -5515 5795
rect -5535 5570 -5515 5775
rect -4925 5705 -4905 5900
rect -5535 5550 -5440 5570
rect -5075 5550 -4945 5570
rect -5660 5500 -5480 5520
rect -5660 5225 -5525 5245
rect -5545 5065 -5525 5225
rect -5500 5220 -5480 5500
rect -4965 5240 -4945 5550
rect -4965 5220 -4915 5240
rect -5500 5200 -5430 5220
rect -5070 5200 -4985 5220
rect -5005 5195 -4985 5200
rect -5005 5175 -4955 5195
rect -5545 5045 -5475 5065
rect -5660 4950 -5525 4970
rect -5660 4675 -5640 4695
rect -5545 4520 -5525 4950
rect -5495 4870 -5475 5045
rect -5495 4850 -5435 4870
rect -5090 4850 -4995 4870
rect -5545 4500 -5415 4520
rect -5075 4500 -5035 4520
rect -5660 4400 -5640 4420
rect -5660 4125 -5640 4145
rect -5660 3850 -5640 3870
rect -5660 3575 -5640 3595
rect -5055 3540 -5035 4500
rect -5015 3585 -4995 4850
rect -4975 3630 -4955 5175
rect -4935 4105 -4915 5220
rect -4975 3610 -4890 3630
rect -5015 3565 -4945 3585
rect -5055 3520 -4990 3540
rect -5660 3300 -5640 3320
rect -5660 3025 -5640 3045
rect -5660 2750 -5640 2770
rect -5765 2130 -5610 2145
rect -5765 2100 -5750 2130
rect -5630 2100 -5610 2130
rect -7290 1995 -6230 2035
rect -5765 1980 -5610 2100
rect -5765 1950 -5745 1980
rect -5625 1950 -5610 1980
rect -5010 1990 -4990 3520
rect -4965 2035 -4945 3565
rect -4910 2540 -4890 3610
rect -4925 2500 -4890 2540
rect -4965 2015 -4865 2035
rect -5010 1970 -4945 1990
rect -5765 1935 -5610 1950
rect -7290 990 -7180 1025
rect -7275 900 -7235 910
rect -7275 850 -7265 900
rect -7245 850 -7235 900
rect -7275 765 -7235 850
rect -5190 745 -5085 780
rect -5125 680 -5085 745
rect -4965 750 -4945 1970
rect -4885 1400 -4865 2015
rect -4925 1350 -4865 1400
rect -4965 720 -4810 750
rect -5125 630 -5115 680
rect -5095 630 -5085 680
rect -5125 620 -5085 630
rect 2745 680 2785 790
rect 2745 630 2755 680
rect 2775 630 2785 680
rect 2745 620 2785 630
<< viali >>
rect -5980 7030 -5960 7080
rect -5980 6905 -5920 6925
rect -5750 2100 -5630 2130
rect -5745 1950 -5625 1980
rect -7265 850 -7245 900
rect -5115 630 -5095 680
rect 2755 630 2775 680
<< metal1 >>
rect -4545 8735 -4395 8775
rect -7290 8115 -7065 8715
rect -4995 8690 -4530 8715
rect -4995 8115 -4870 8690
rect -4660 8675 -4530 8690
rect -4660 8670 -4595 8675
rect -7290 7425 -7065 8015
rect -7290 6875 -6690 6920
rect -6730 6835 -6690 6875
rect -6645 6845 -6185 7480
rect -4910 7250 -4870 8115
rect -5990 7205 -4870 7250
rect -5990 7080 -5950 7205
rect -5990 7030 -5980 7080
rect -5960 7030 -5950 7080
rect -5990 7020 -5950 7030
rect -5465 6975 -5050 7205
rect -5990 6925 -5910 6935
rect -5990 6905 -5980 6925
rect -5920 6905 -5910 6925
rect -5990 6880 -5910 6905
rect -6130 6830 -5660 6880
rect -5545 6865 -5050 6975
rect -5545 6795 -5365 6865
rect -5545 6535 -5490 6795
rect -5065 6640 -4785 6730
rect -5545 6445 -5385 6535
rect -5545 6185 -5490 6445
rect -5070 6290 -4790 6380
rect -5545 6095 -5440 6185
rect -5545 5835 -5490 6095
rect -5065 5940 -4785 6030
rect -5545 5745 -5440 5835
rect -5545 5485 -5490 5745
rect -5065 5590 -4785 5680
rect -5545 5395 -5440 5485
rect -5545 5135 -5490 5395
rect -5065 5240 -4785 5330
rect -5545 5045 -5440 5135
rect -5545 4785 -5490 5045
rect -5065 4890 -4785 4980
rect -5545 4695 -5440 4785
rect -5065 4540 -4785 4630
rect -6640 2275 -6185 2430
rect -5660 2350 -5610 2380
rect -6640 2130 -4810 2275
rect -6640 2100 -5750 2130
rect -5630 2100 -4810 2130
rect -6640 2095 -4810 2100
rect -5765 2085 -4810 2095
rect -7275 2020 -5015 2060
rect -7275 900 -7235 2020
rect -5765 1980 -5475 2000
rect -5765 1950 -5745 1980
rect -5625 1950 -5475 1980
rect -5765 1915 -5475 1950
rect -7275 850 -7265 900
rect -7245 850 -7235 900
rect -7275 830 -7235 850
rect -5125 680 -5085 690
rect -5125 630 -5115 680
rect -5095 630 -5085 680
rect -5125 550 -5085 630
rect -5060 605 -5015 2020
rect 2810 785 2905 830
rect 2745 680 2785 690
rect 2745 630 2755 680
rect 2775 630 2785 680
rect 2745 605 2785 630
rect -5060 565 2785 605
rect 2860 550 2905 785
rect -5125 505 2905 550
use dac  dac_0 ~/VLSI_Sine_Gen/layout/dac
timestamp 1702787255
transform 1 0 -4510 0 1 7245
box -415 -6625 7355 1590
use filter  filter_0 ~/VLSI_Sine_Gen/layout/filter
timestamp 1702883810
transform 1 0 -6820 0 1 135
box -420 455 1685 1890
use inverter  inverter_0 ~/VLSI_Sine_Gen/layout/dac
timestamp 1693780072
transform 1 0 -5020 0 1 4625
box -240 -145 -30 185
use inverter  inverter_1
timestamp 1693780072
transform 1 0 -5225 0 1 6725
box -240 -145 -30 185
use inverter  inverter_2
timestamp 1693780072
transform 1 0 -5225 0 1 4625
box -240 -145 -30 185
use inverter  inverter_3
timestamp 1693780072
transform 1 0 -5225 0 1 6375
box -240 -145 -30 185
use inverter  inverter_4
timestamp 1693780072
transform 1 0 -5225 0 1 6025
box -240 -145 -30 185
use inverter  inverter_5
timestamp 1693780072
transform 1 0 -5020 0 1 6725
box -240 -145 -30 185
use inverter  inverter_6
timestamp 1693780072
transform 1 0 -5020 0 1 6375
box -240 -145 -30 185
use inverter  inverter_7
timestamp 1693780072
transform 1 0 -5020 0 1 6025
box -240 -145 -30 185
use inverter  inverter_8
timestamp 1693780072
transform 1 0 -5225 0 1 5675
box -240 -145 -30 185
use inverter  inverter_9
timestamp 1693780072
transform 1 0 -5225 0 1 5325
box -240 -145 -30 185
use inverter  inverter_10
timestamp 1693780072
transform 1 0 -5225 0 1 4975
box -240 -145 -30 185
use inverter  inverter_11
timestamp 1693780072
transform 1 0 -5020 0 1 5675
box -240 -145 -30 185
use inverter  inverter_12
timestamp 1693780072
transform 1 0 -5020 0 1 5325
box -240 -145 -30 185
use inverter  inverter_13
timestamp 1693780072
transform 1 0 -5020 0 1 4975
box -240 -145 -30 185
use register16  register16_0 ~/VLSI_Sine_Gen/layout/shift_register
timestamp 1702679440
transform 0 1 -6715 -1 0 6885
box -90 -15 4570 1140
use v_gen  v_gen_0 ~/VLSI_Sine_Gen/layout/v_gen
timestamp 1702787459
transform 1 0 -7075 0 1 7375
box -35 -10 2120 1435
<< labels >>
rlabel metal1 -5610 2365 -5610 2365 3 Vff16
port 22 e
rlabel locali -5640 4685 -5640 4685 3 Vff8
port 14 e
rlabel locali -5640 4410 -5640 4410 3 Vff9
port 15 e
rlabel locali -5640 4135 -5640 4135 3 Vff10
port 16 e
rlabel locali -5640 3860 -5640 3860 3 Vff11
port 17 e
rlabel locali -5640 3585 -5640 3585 3 Vff12
port 18 e
rlabel locali -5640 3310 -5640 3310 3 Vff13
port 19 e
rlabel locali -5640 3035 -5640 3035 3 Vff14
port 20 e
rlabel locali -5640 2760 -5640 2760 3 Vff15
port 21 e
rlabel locali -5575 6610 -5575 6610 3 Vphi1
port 7 e
rlabel locali -5575 6335 -5575 6335 3 Vphi2
port 8 e
rlabel locali -5575 6060 -5575 6060 3 Vphi3
port 9 e
rlabel locali -5575 5785 -5575 5785 3 Vphi4
port 10 e
rlabel locali -5575 5510 -5575 5510 3 Vphi5
port 11 e
rlabel locali -5575 5235 -5575 5235 3 Vphi6
port 12 e
rlabel locali -5575 4960 -5575 4960 3 Vphi7
port 13 e
rlabel locali -7290 2015 -7290 2015 7 Voutn
port 6 w
rlabel locali -7290 1005 -7290 1005 7 Voutp
port 5 w
rlabel metal1 -7290 6895 -7290 6895 1 CLK
port 2 n
rlabel metal1 -7290 8415 -7290 8415 7 VP
port 3 w
rlabel metal1 -7290 7720 -7290 7720 7 VN
port 4 w
rlabel locali -7290 7375 -7290 7375 7 Vb
port 1 w
<< end >>
