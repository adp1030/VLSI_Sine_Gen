magic
tech sky130A
timestamp 1702636620
<< nwell >>
rect 4835 105 4950 1460
rect 5635 -1495 5755 -140
rect 5635 -4700 5765 -3345
rect 4835 -6305 4975 -4950
<< poly >>
rect 5975 1575 6025 1585
rect -15 1560 6025 1575
rect -15 -25 0 1560
rect 270 1430 320 1560
rect 370 1520 420 1530
rect 370 1500 380 1520
rect 410 1500 420 1520
rect 370 1430 420 1500
rect 1070 1430 1120 1560
rect 1170 1520 1220 1530
rect 1170 1500 1180 1520
rect 1210 1500 1220 1520
rect 1170 1435 1220 1500
rect 1870 1430 1920 1560
rect 1970 1520 2020 1530
rect 1970 1500 1980 1520
rect 2010 1500 2020 1520
rect 1970 1435 2020 1500
rect 2670 1430 2720 1560
rect 2770 1520 2820 1530
rect 2770 1500 2780 1520
rect 2810 1500 2820 1520
rect 2770 1435 2820 1500
rect 3470 1430 3520 1560
rect 3570 1520 3620 1530
rect 3570 1500 3580 1520
rect 3610 1500 3620 1520
rect 3570 1435 3620 1500
rect 4270 1430 4320 1560
rect 4370 1520 4420 1530
rect 4370 1500 4380 1520
rect 4410 1500 4420 1520
rect 4370 1435 4420 1500
rect 5175 1430 5225 1560
rect 5275 1520 5325 1530
rect 5275 1500 5285 1520
rect 5315 1500 5325 1520
rect 5275 1435 5325 1500
rect 5975 1430 6025 1560
rect 6075 1530 6125 1585
rect 6075 1520 6655 1530
rect 6075 1500 6085 1520
rect 6115 1515 6655 1520
rect 6115 1500 6125 1515
rect 6075 1435 6125 1500
rect -15 -40 6025 -25
rect -15 -1625 0 -40
rect 270 -165 320 -40
rect 990 -75 1040 -65
rect 990 -80 1000 -75
rect 370 -95 1000 -80
rect 1030 -95 1040 -75
rect 370 -100 1040 -95
rect 370 -165 420 -100
rect 990 -105 1040 -100
rect 1070 -165 1120 -40
rect 1170 -75 1220 -65
rect 1170 -95 1180 -75
rect 1210 -80 1220 -75
rect 1790 -75 1840 -65
rect 1790 -80 1800 -75
rect 1210 -95 1800 -80
rect 1830 -95 1840 -75
rect 1170 -100 1840 -95
rect 1170 -165 1220 -100
rect 1790 -105 1840 -100
rect 1870 -165 1920 -40
rect 1970 -75 2020 -65
rect 1970 -95 1980 -75
rect 2010 -80 2020 -75
rect 2590 -75 2640 -65
rect 2590 -80 2600 -75
rect 2010 -95 2600 -80
rect 2630 -95 2640 -75
rect 1970 -100 2640 -95
rect 1970 -165 2020 -100
rect 2590 -105 2640 -100
rect 2670 -165 2720 -40
rect 2770 -75 2820 -65
rect 2770 -95 2780 -75
rect 2810 -80 2820 -75
rect 3390 -75 3440 -65
rect 3390 -80 3400 -75
rect 2810 -95 3400 -80
rect 3430 -95 3440 -75
rect 2770 -100 3440 -95
rect 2770 -165 2820 -100
rect 3390 -105 3440 -100
rect 3470 -165 3520 -40
rect 3570 -75 3620 -65
rect 3570 -95 3580 -75
rect 3610 -80 3620 -75
rect 4190 -75 4240 -65
rect 4190 -80 4200 -75
rect 3610 -95 4200 -80
rect 4230 -95 4240 -75
rect 3570 -100 4240 -95
rect 3570 -165 3620 -100
rect 4190 -105 4240 -100
rect 4270 -165 4320 -40
rect 4370 -75 4420 -65
rect 4370 -95 4380 -75
rect 4410 -80 4420 -75
rect 4990 -75 5040 -65
rect 4990 -80 5000 -75
rect 4410 -95 5000 -80
rect 5030 -95 5040 -75
rect 4370 -100 5040 -95
rect 4370 -165 4420 -100
rect 4990 -105 5040 -100
rect 5070 -165 5120 -40
rect 5170 -75 5220 -65
rect 5170 -95 5180 -75
rect 5210 -80 5220 -75
rect 5895 -75 5945 -65
rect 5895 -80 5905 -75
rect 5210 -95 5905 -80
rect 5935 -95 5945 -75
rect 5170 -100 5945 -95
rect 5170 -165 5220 -100
rect 5895 -105 5945 -100
rect 5975 -165 6025 -40
rect 6075 -75 6125 -65
rect 6075 -95 6085 -75
rect 6115 -80 6125 -75
rect 6640 -80 6655 1515
rect 6115 -95 6655 -80
rect 6075 -100 6655 -95
rect 6075 -165 6125 -100
rect -15 -1640 5920 -1625
rect -15 -3225 0 -1640
rect 270 -1765 320 -1640
rect 370 -1680 420 -1665
rect 990 -1675 1040 -1665
rect 990 -1680 1000 -1675
rect 370 -1695 1000 -1680
rect 1030 -1695 1040 -1675
rect 370 -1700 1040 -1695
rect 370 -1765 420 -1700
rect 990 -1705 1040 -1700
rect 1070 -1765 1120 -1640
rect 1170 -1675 1220 -1665
rect 1170 -1695 1180 -1675
rect 1210 -1680 1220 -1675
rect 1790 -1675 1840 -1665
rect 1790 -1680 1800 -1675
rect 1210 -1695 1800 -1680
rect 1830 -1695 1840 -1675
rect 1170 -1700 1840 -1695
rect 1170 -1765 1220 -1700
rect 1790 -1705 1840 -1700
rect 1870 -1765 1920 -1640
rect 1970 -1675 2020 -1665
rect 1970 -1695 1980 -1675
rect 2010 -1680 2020 -1675
rect 2590 -1675 2640 -1665
rect 2590 -1680 2600 -1675
rect 2010 -1695 2600 -1680
rect 2630 -1695 2640 -1675
rect 1970 -1700 2640 -1695
rect 1970 -1770 2020 -1700
rect 2590 -1705 2640 -1700
rect 2670 -1765 2720 -1640
rect 2770 -1675 2820 -1665
rect 2770 -1695 2780 -1675
rect 2810 -1680 2820 -1675
rect 3390 -1675 3440 -1665
rect 3390 -1680 3400 -1675
rect 2810 -1695 3400 -1680
rect 3430 -1695 3440 -1675
rect 2770 -1700 3440 -1695
rect 2770 -1765 2820 -1700
rect 3390 -1705 3440 -1700
rect 3470 -1765 3520 -1640
rect 3570 -1675 3620 -1665
rect 3570 -1695 3580 -1675
rect 3610 -1680 3620 -1675
rect 4190 -1675 4240 -1665
rect 4190 -1680 4200 -1675
rect 3610 -1695 4200 -1680
rect 4230 -1695 4240 -1675
rect 3570 -1700 4240 -1695
rect 3570 -1765 3620 -1700
rect 4190 -1705 4240 -1700
rect 4270 -1765 4320 -1640
rect 4370 -1675 4420 -1665
rect 4370 -1695 4380 -1675
rect 4410 -1680 4420 -1675
rect 4990 -1675 5040 -1665
rect 4990 -1680 5000 -1675
rect 4410 -1695 5000 -1680
rect 5030 -1695 5040 -1675
rect 4370 -1700 5040 -1695
rect 4370 -1765 4420 -1700
rect 4990 -1705 5040 -1700
rect 5070 -1765 5120 -1640
rect 5170 -1675 5220 -1665
rect 5170 -1695 5180 -1675
rect 5210 -1680 5220 -1675
rect 5790 -1675 5840 -1665
rect 5790 -1680 5800 -1675
rect 5210 -1695 5800 -1680
rect 5830 -1695 5840 -1675
rect 5170 -1700 5840 -1695
rect 5170 -1765 5220 -1700
rect 5790 -1705 5840 -1700
rect 5870 -1765 5920 -1640
rect 5970 -1675 6020 -1665
rect 5970 -1695 5980 -1675
rect 6010 -1680 6020 -1675
rect 6640 -1680 6655 -100
rect 6010 -1695 6655 -1680
rect 5970 -1700 6655 -1695
rect 5970 -1765 6020 -1700
rect -15 -3240 6025 -3225
rect -15 -4830 0 -3240
rect 270 -3370 320 -3240
rect 370 -3280 420 -3265
rect 990 -3275 1040 -3265
rect 990 -3280 1000 -3275
rect 370 -3295 1000 -3280
rect 1030 -3295 1040 -3275
rect 370 -3300 1040 -3295
rect 370 -3370 420 -3300
rect 990 -3305 1040 -3300
rect 1070 -3370 1120 -3240
rect 1170 -3275 1220 -3265
rect 1170 -3295 1180 -3275
rect 1210 -3280 1220 -3275
rect 1790 -3275 1840 -3265
rect 1790 -3280 1800 -3275
rect 1210 -3295 1800 -3280
rect 1830 -3295 1840 -3275
rect 1170 -3300 1840 -3295
rect 1170 -3370 1220 -3300
rect 1790 -3305 1840 -3300
rect 1870 -3375 1920 -3240
rect 1970 -3275 2020 -3265
rect 1970 -3295 1980 -3275
rect 2010 -3280 2020 -3275
rect 2590 -3275 2640 -3265
rect 2590 -3280 2600 -3275
rect 2010 -3295 2600 -3280
rect 2630 -3295 2640 -3275
rect 1970 -3300 2640 -3295
rect 1970 -3370 2020 -3300
rect 2590 -3305 2640 -3300
rect 2670 -3370 2720 -3240
rect 2770 -3275 2820 -3265
rect 2770 -3295 2780 -3275
rect 2810 -3280 2820 -3275
rect 3390 -3275 3440 -3265
rect 3390 -3280 3400 -3275
rect 2810 -3295 3400 -3280
rect 3430 -3295 3440 -3275
rect 2770 -3300 3440 -3295
rect 2770 -3370 2820 -3300
rect 3390 -3305 3440 -3300
rect 3470 -3370 3520 -3240
rect 3570 -3275 3620 -3265
rect 3570 -3295 3580 -3275
rect 3610 -3280 3620 -3275
rect 4190 -3275 4240 -3265
rect 4190 -3280 4200 -3275
rect 3610 -3295 4200 -3280
rect 4230 -3295 4240 -3275
rect 3570 -3300 4240 -3295
rect 3570 -3370 3620 -3300
rect 4190 -3305 4240 -3300
rect 4270 -3370 4320 -3240
rect 4370 -3275 4420 -3265
rect 4370 -3295 4380 -3275
rect 4410 -3280 4420 -3275
rect 4990 -3275 5040 -3265
rect 4990 -3280 5000 -3275
rect 4410 -3295 5000 -3280
rect 5030 -3295 5040 -3275
rect 4370 -3300 5040 -3295
rect 4370 -3370 4420 -3300
rect 4990 -3305 5040 -3300
rect 5070 -3370 5120 -3240
rect 5170 -3275 5220 -3265
rect 5170 -3295 5180 -3275
rect 5210 -3280 5220 -3275
rect 5895 -3275 5945 -3265
rect 5895 -3280 5905 -3275
rect 5210 -3295 5905 -3280
rect 5935 -3295 5945 -3275
rect 5170 -3300 5945 -3295
rect 5170 -3370 5220 -3300
rect 5895 -3305 5945 -3300
rect 5975 -3370 6025 -3240
rect 6075 -3275 6125 -3265
rect 6075 -3295 6085 -3275
rect 6115 -3280 6125 -3275
rect 6640 -3280 6655 -1700
rect 6115 -3295 6655 -3280
rect 6075 -3300 6655 -3295
rect 6075 -3370 6125 -3300
rect -15 -4845 6025 -4830
rect 270 -4975 320 -4845
rect 370 -4885 420 -4870
rect 990 -4880 1040 -4870
rect 990 -4885 1000 -4880
rect 370 -4900 1000 -4885
rect 1030 -4900 1040 -4880
rect 370 -4905 1040 -4900
rect 370 -4975 420 -4905
rect 990 -4910 1040 -4905
rect 1070 -4975 1120 -4845
rect 1170 -4880 1220 -4870
rect 1170 -4900 1180 -4880
rect 1210 -4885 1220 -4880
rect 1790 -4880 1840 -4870
rect 1790 -4885 1800 -4880
rect 1210 -4900 1800 -4885
rect 1830 -4900 1840 -4880
rect 1170 -4905 1840 -4900
rect 1170 -4975 1220 -4905
rect 1790 -4910 1840 -4905
rect 1870 -4975 1920 -4845
rect 1970 -4880 2020 -4870
rect 1970 -4900 1980 -4880
rect 2010 -4885 2020 -4880
rect 2590 -4880 2640 -4870
rect 2590 -4885 2600 -4880
rect 2010 -4900 2600 -4885
rect 2630 -4900 2640 -4880
rect 1970 -4905 2640 -4900
rect 1970 -4975 2020 -4905
rect 2590 -4910 2640 -4905
rect 2670 -4975 2720 -4845
rect 2770 -4880 2820 -4870
rect 2770 -4900 2780 -4880
rect 2810 -4885 2820 -4880
rect 3390 -4880 3440 -4870
rect 3390 -4885 3400 -4880
rect 2810 -4900 3400 -4885
rect 3430 -4900 3440 -4880
rect 2770 -4905 3440 -4900
rect 2770 -4975 2820 -4905
rect 3390 -4910 3440 -4905
rect 3470 -4975 3520 -4845
rect 3570 -4880 3620 -4870
rect 3570 -4900 3580 -4880
rect 3610 -4885 3620 -4880
rect 4190 -4880 4240 -4870
rect 4190 -4885 4200 -4880
rect 3610 -4900 4200 -4885
rect 4230 -4900 4240 -4880
rect 3570 -4905 4240 -4900
rect 3570 -4975 3620 -4905
rect 4190 -4910 4240 -4905
rect 4270 -4975 4320 -4845
rect 4370 -4880 4420 -4870
rect 4370 -4900 4380 -4880
rect 4410 -4885 4420 -4880
rect 5095 -4880 5145 -4870
rect 5095 -4885 5105 -4880
rect 4410 -4900 5105 -4885
rect 5135 -4900 5145 -4880
rect 4370 -4905 5145 -4900
rect 4370 -4975 4420 -4905
rect 5095 -4910 5145 -4905
rect 5175 -4975 5225 -4845
rect 5275 -4880 5325 -4870
rect 5275 -4900 5285 -4880
rect 5315 -4885 5325 -4880
rect 5895 -4880 5945 -4870
rect 5895 -4885 5905 -4880
rect 5315 -4900 5905 -4885
rect 5935 -4900 5945 -4880
rect 5275 -4905 5945 -4900
rect 5275 -4975 5325 -4905
rect 5895 -4910 5945 -4905
rect 5975 -4975 6025 -4845
rect 6075 -4880 6125 -4870
rect 6075 -4900 6085 -4880
rect 6115 -4885 6125 -4880
rect 6640 -4885 6655 -3300
rect 6115 -4900 6655 -4885
rect 6075 -4905 6655 -4900
rect 6075 -4975 6125 -4905
<< polycont >>
rect 380 1500 410 1520
rect 1180 1500 1210 1520
rect 1980 1500 2010 1520
rect 2780 1500 2810 1520
rect 3580 1500 3610 1520
rect 4380 1500 4410 1520
rect 5285 1500 5315 1520
rect 6085 1500 6115 1520
rect 1000 -95 1030 -75
rect 1180 -95 1210 -75
rect 1800 -95 1830 -75
rect 1980 -95 2010 -75
rect 2600 -95 2630 -75
rect 2780 -95 2810 -75
rect 3400 -95 3430 -75
rect 3580 -95 3610 -75
rect 4200 -95 4230 -75
rect 4380 -95 4410 -75
rect 5000 -95 5030 -75
rect 5180 -95 5210 -75
rect 5905 -95 5935 -75
rect 6085 -95 6115 -75
rect 1000 -1695 1030 -1675
rect 1180 -1695 1210 -1675
rect 1800 -1695 1830 -1675
rect 1980 -1695 2010 -1675
rect 2600 -1695 2630 -1675
rect 2780 -1695 2810 -1675
rect 3400 -1695 3430 -1675
rect 3580 -1695 3610 -1675
rect 4200 -1695 4230 -1675
rect 4380 -1695 4410 -1675
rect 5000 -1695 5030 -1675
rect 5180 -1695 5210 -1675
rect 5800 -1695 5830 -1675
rect 5980 -1695 6010 -1675
rect 1000 -3295 1030 -3275
rect 1180 -3295 1210 -3275
rect 1800 -3295 1830 -3275
rect 1980 -3295 2010 -3275
rect 2600 -3295 2630 -3275
rect 2780 -3295 2810 -3275
rect 3400 -3295 3430 -3275
rect 3580 -3295 3610 -3275
rect 4200 -3295 4230 -3275
rect 4380 -3295 4410 -3275
rect 5000 -3295 5030 -3275
rect 5180 -3295 5210 -3275
rect 5905 -3295 5935 -3275
rect 6085 -3295 6115 -3275
rect 1000 -4900 1030 -4880
rect 1180 -4900 1210 -4880
rect 1800 -4900 1830 -4880
rect 1980 -4900 2010 -4880
rect 2600 -4900 2630 -4880
rect 2780 -4900 2810 -4880
rect 3400 -4900 3430 -4880
rect 3580 -4900 3610 -4880
rect 4200 -4900 4230 -4880
rect 4380 -4900 4410 -4880
rect 5105 -4900 5135 -4880
rect 5285 -4900 5315 -4880
rect 5905 -4900 5935 -4880
rect 6085 -4900 6115 -4880
<< locali >>
rect 370 1520 6125 1530
rect 370 1500 380 1520
rect 410 1500 1180 1520
rect 1210 1500 1980 1520
rect 2010 1500 2780 1520
rect 2810 1500 3580 1520
rect 3610 1500 4380 1520
rect 4410 1500 5285 1520
rect 5315 1500 6085 1520
rect 6115 1500 6125 1520
rect 370 1495 6125 1500
rect 370 1490 420 1495
rect 1170 1490 1220 1495
rect 1970 1490 2020 1495
rect 2770 1490 2820 1495
rect 3570 1490 3620 1495
rect 4370 1490 4420 1495
rect 5275 1490 5325 1495
rect 6075 1490 6125 1495
rect 6625 175 6665 185
rect 6625 125 6635 175
rect 6655 125 6665 175
rect 6625 45 6665 125
rect 225 -65 260 45
rect 430 -10 460 45
rect 430 -20 500 -10
rect 430 -40 440 -20
rect 490 -40 500 -20
rect 430 -50 500 -40
rect 920 -15 1060 20
rect 1230 -10 1260 45
rect 1825 20 1860 45
rect 920 -65 955 -15
rect 1230 -20 1300 -10
rect 1230 -40 1240 -20
rect 1290 -40 1300 -20
rect 1230 -50 1300 -40
rect 1720 -15 1860 20
rect 2030 -10 2060 45
rect 2625 20 2660 45
rect 1720 -65 1755 -15
rect 2030 -20 2100 -10
rect 2030 -40 2040 -20
rect 2090 -40 2100 -20
rect 2030 -50 2100 -40
rect 2520 -15 2660 20
rect 2830 -10 2860 45
rect 3425 20 3460 45
rect 2520 -65 2555 -15
rect 2830 -20 2900 -10
rect 2830 -40 2840 -20
rect 2890 -40 2900 -20
rect 2830 -50 2900 -40
rect 3320 -15 3460 20
rect 3630 -10 3660 45
rect 4225 20 4260 45
rect 3320 -65 3355 -15
rect 3630 -20 3700 -10
rect 3630 -40 3640 -20
rect 3690 -40 3700 -20
rect 3630 -50 3700 -40
rect 4120 -15 4260 20
rect 4430 -10 4460 45
rect 5130 20 5165 45
rect 4120 -65 4155 -15
rect 4430 -20 4500 -10
rect 4430 -40 4440 -20
rect 4490 -40 4500 -20
rect 4430 -50 4500 -40
rect 4920 -15 5165 20
rect 5335 -10 5365 45
rect 5930 20 5965 45
rect 4920 -65 4955 -15
rect 5235 -20 5365 -10
rect 5235 -40 5245 -20
rect 5295 -35 5365 -20
rect 5825 -15 5965 20
rect 6135 -10 6165 45
rect 6595 40 6665 45
rect 6595 20 6605 40
rect 6655 20 6665 40
rect 6595 10 6665 20
rect 5295 -40 5305 -35
rect 5235 -50 5305 -40
rect 5825 -65 5860 -15
rect 6135 -20 6205 -10
rect 6135 -40 6145 -20
rect 6195 -40 6205 -20
rect 6135 -50 6205 -40
rect 6595 -20 6885 -10
rect 6595 -40 6605 -20
rect 6655 -40 6825 -20
rect 6875 -40 6885 -20
rect 6595 -50 6885 -40
rect 225 -75 295 -65
rect 225 -95 235 -75
rect 285 -95 295 -75
rect 225 -105 295 -95
rect 885 -75 955 -65
rect 885 -95 895 -75
rect 945 -95 955 -75
rect 885 -105 955 -95
rect 990 -75 1220 -65
rect 990 -95 1000 -75
rect 1030 -95 1180 -75
rect 1210 -95 1220 -75
rect 990 -105 1220 -95
rect 1685 -75 1755 -65
rect 1685 -95 1695 -75
rect 1745 -95 1755 -75
rect 1685 -105 1755 -95
rect 1790 -75 2020 -65
rect 1790 -95 1800 -75
rect 1830 -95 1980 -75
rect 2010 -95 2020 -75
rect 1790 -105 2020 -95
rect 2485 -75 2555 -65
rect 2485 -95 2495 -75
rect 2545 -95 2555 -75
rect 2485 -105 2555 -95
rect 2590 -75 2820 -65
rect 2590 -95 2600 -75
rect 2630 -95 2780 -75
rect 2810 -95 2820 -75
rect 2590 -105 2820 -95
rect 3285 -75 3355 -65
rect 3285 -95 3295 -75
rect 3345 -95 3355 -75
rect 3285 -105 3355 -95
rect 3390 -75 3620 -65
rect 3390 -95 3400 -75
rect 3430 -95 3580 -75
rect 3610 -95 3620 -75
rect 3390 -105 3620 -95
rect 4085 -75 4155 -65
rect 4085 -95 4095 -75
rect 4145 -95 4155 -75
rect 4085 -105 4155 -95
rect 4190 -75 4420 -65
rect 4190 -95 4200 -75
rect 4230 -95 4380 -75
rect 4410 -95 4420 -75
rect 4190 -105 4420 -95
rect 4885 -75 4955 -65
rect 4885 -95 4895 -75
rect 4945 -95 4955 -75
rect 4885 -105 4955 -95
rect 4990 -75 5220 -65
rect 4990 -95 5000 -75
rect 5030 -95 5180 -75
rect 5210 -95 5220 -75
rect 4990 -105 5220 -95
rect 5790 -75 5860 -65
rect 5790 -95 5800 -75
rect 5850 -95 5860 -75
rect 5790 -105 5860 -95
rect 5895 -75 6125 -65
rect 5895 -95 5905 -75
rect 5935 -95 6085 -75
rect 6115 -95 6125 -75
rect 5895 -105 6125 -95
rect 6625 -85 6665 -75
rect 6625 -135 6635 -85
rect 6655 -105 6665 -85
rect 6655 -115 6830 -105
rect 6655 -135 6800 -115
rect 6625 -145 6800 -135
rect 6790 -165 6800 -145
rect 6820 -165 6830 -115
rect 6790 -175 6830 -165
rect 6735 -1445 6775 -1435
rect 6735 -1470 6745 -1445
rect 6625 -1480 6745 -1470
rect 6625 -1530 6635 -1480
rect 6655 -1495 6745 -1480
rect 6765 -1495 6775 -1445
rect 6655 -1505 6775 -1495
rect 6655 -1530 6665 -1505
rect 6625 -1540 6665 -1530
rect 6790 -1535 6830 -1525
rect 225 -1665 260 -1555
rect 430 -1610 460 -1555
rect 430 -1620 500 -1610
rect 430 -1640 440 -1620
rect 490 -1640 500 -1620
rect 430 -1650 500 -1640
rect 920 -1615 1060 -1580
rect 1230 -1610 1260 -1555
rect 920 -1665 955 -1615
rect 1230 -1620 1300 -1610
rect 1230 -1640 1240 -1620
rect 1290 -1640 1300 -1620
rect 1230 -1650 1300 -1640
rect 1720 -1615 1860 -1580
rect 2030 -1610 2060 -1555
rect 1720 -1665 1755 -1615
rect 2030 -1620 2100 -1610
rect 2030 -1640 2040 -1620
rect 2090 -1640 2100 -1620
rect 2030 -1650 2100 -1640
rect 2520 -1615 2660 -1580
rect 2830 -1610 2860 -1555
rect 2520 -1665 2555 -1615
rect 2830 -1620 2900 -1610
rect 2830 -1640 2840 -1620
rect 2890 -1640 2900 -1620
rect 2830 -1650 2900 -1640
rect 3320 -1615 3460 -1580
rect 3630 -1610 3660 -1555
rect 3320 -1665 3355 -1615
rect 3630 -1620 3700 -1610
rect 3630 -1640 3640 -1620
rect 3690 -1640 3700 -1620
rect 3630 -1650 3700 -1640
rect 4120 -1615 4260 -1580
rect 4430 -1610 4460 -1555
rect 4120 -1665 4155 -1615
rect 4430 -1620 4500 -1610
rect 4430 -1640 4440 -1620
rect 4490 -1640 4500 -1620
rect 4430 -1650 4500 -1640
rect 4920 -1615 5060 -1580
rect 5230 -1610 5260 -1555
rect 4920 -1665 4955 -1615
rect 5230 -1620 5300 -1610
rect 5230 -1640 5240 -1620
rect 5290 -1640 5300 -1620
rect 5230 -1650 5300 -1640
rect 5720 -1615 5965 -1580
rect 6135 -1610 6165 -1550
rect 5720 -1665 5755 -1615
rect 6035 -1620 6165 -1610
rect 6035 -1640 6045 -1620
rect 6095 -1640 6165 -1620
rect 6035 -1650 6165 -1640
rect 6790 -1585 6800 -1535
rect 6820 -1585 6830 -1535
rect 6790 -1665 6830 -1585
rect 225 -1675 295 -1665
rect 225 -1695 235 -1675
rect 285 -1695 295 -1675
rect 225 -1705 295 -1695
rect 885 -1675 955 -1665
rect 885 -1695 895 -1675
rect 945 -1695 955 -1675
rect 885 -1705 955 -1695
rect 990 -1675 1220 -1665
rect 990 -1695 1000 -1675
rect 1030 -1695 1180 -1675
rect 1210 -1695 1220 -1675
rect 990 -1705 1220 -1695
rect 1685 -1675 1755 -1665
rect 1685 -1695 1695 -1675
rect 1745 -1695 1755 -1675
rect 1685 -1705 1755 -1695
rect 1790 -1675 2020 -1665
rect 1790 -1695 1800 -1675
rect 1830 -1695 1980 -1675
rect 2010 -1695 2020 -1675
rect 1790 -1705 2020 -1695
rect 2485 -1675 2555 -1665
rect 2485 -1695 2495 -1675
rect 2545 -1695 2555 -1675
rect 2485 -1705 2555 -1695
rect 2590 -1675 2820 -1665
rect 2590 -1695 2600 -1675
rect 2630 -1695 2780 -1675
rect 2810 -1695 2820 -1675
rect 2590 -1705 2820 -1695
rect 3285 -1675 3355 -1665
rect 3285 -1695 3295 -1675
rect 3345 -1695 3355 -1675
rect 3285 -1705 3355 -1695
rect 3390 -1675 3620 -1665
rect 3390 -1695 3400 -1675
rect 3430 -1695 3580 -1675
rect 3610 -1695 3620 -1675
rect 3390 -1705 3620 -1695
rect 4085 -1675 4155 -1665
rect 4085 -1695 4095 -1675
rect 4145 -1695 4155 -1675
rect 4085 -1705 4155 -1695
rect 4190 -1675 4420 -1665
rect 4190 -1695 4200 -1675
rect 4230 -1695 4380 -1675
rect 4410 -1695 4420 -1675
rect 4190 -1705 4420 -1695
rect 4885 -1675 4955 -1665
rect 4885 -1695 4895 -1675
rect 4945 -1695 4955 -1675
rect 4885 -1705 4955 -1695
rect 4990 -1675 5220 -1665
rect 4990 -1695 5000 -1675
rect 5030 -1695 5180 -1675
rect 5210 -1695 5220 -1675
rect 4990 -1705 5220 -1695
rect 5685 -1675 5755 -1665
rect 5685 -1695 5695 -1675
rect 5745 -1695 5755 -1675
rect 5685 -1705 5755 -1695
rect 5790 -1675 6020 -1665
rect 5790 -1695 5800 -1675
rect 5830 -1695 5980 -1675
rect 6010 -1695 6020 -1675
rect 5790 -1705 6020 -1695
rect 6760 -1675 6830 -1665
rect 6760 -1695 6770 -1675
rect 6820 -1695 6830 -1675
rect 6760 -1705 6830 -1695
rect 6790 -3135 6830 -3125
rect 225 -3265 260 -3155
rect 430 -3210 460 -3155
rect 430 -3220 500 -3210
rect 430 -3240 440 -3220
rect 490 -3240 500 -3220
rect 430 -3250 500 -3240
rect 920 -3215 1060 -3180
rect 1230 -3210 1260 -3155
rect 920 -3265 955 -3215
rect 1230 -3220 1300 -3210
rect 1230 -3240 1240 -3220
rect 1290 -3240 1300 -3220
rect 1230 -3250 1300 -3240
rect 1720 -3215 1860 -3180
rect 2030 -3210 2060 -3155
rect 1720 -3265 1755 -3215
rect 2030 -3220 2100 -3210
rect 2030 -3240 2040 -3220
rect 2090 -3240 2100 -3220
rect 2030 -3250 2100 -3240
rect 2520 -3215 2660 -3180
rect 2830 -3210 2860 -3155
rect 2520 -3265 2555 -3215
rect 2830 -3220 2900 -3210
rect 2830 -3240 2840 -3220
rect 2890 -3240 2900 -3220
rect 2830 -3250 2900 -3240
rect 3320 -3215 3460 -3180
rect 3630 -3210 3660 -3155
rect 3320 -3265 3355 -3215
rect 3630 -3220 3700 -3210
rect 3630 -3240 3640 -3220
rect 3690 -3240 3700 -3220
rect 3630 -3250 3700 -3240
rect 4120 -3215 4260 -3180
rect 4430 -3210 4460 -3155
rect 4120 -3265 4155 -3215
rect 4430 -3220 4500 -3210
rect 4430 -3240 4440 -3220
rect 4490 -3240 4500 -3220
rect 4430 -3250 4500 -3240
rect 4920 -3215 5060 -3180
rect 5230 -3210 5260 -3155
rect 4920 -3265 4955 -3215
rect 5230 -3220 5300 -3210
rect 5230 -3240 5240 -3220
rect 5290 -3240 5300 -3220
rect 5230 -3250 5300 -3240
rect 5825 -3265 5860 -3175
rect 6030 -3210 6060 -3155
rect 5985 -3220 6060 -3210
rect 5985 -3240 5995 -3220
rect 6045 -3240 6060 -3220
rect 5985 -3250 6060 -3240
rect 6790 -3185 6800 -3135
rect 6820 -3185 6830 -3135
rect 6790 -3265 6830 -3185
rect 225 -3275 295 -3265
rect 225 -3295 235 -3275
rect 285 -3295 295 -3275
rect 225 -3305 295 -3295
rect 885 -3275 955 -3265
rect 885 -3295 895 -3275
rect 945 -3295 955 -3275
rect 885 -3305 955 -3295
rect 990 -3275 1220 -3265
rect 990 -3295 1000 -3275
rect 1030 -3295 1180 -3275
rect 1210 -3295 1220 -3275
rect 990 -3305 1220 -3295
rect 1685 -3275 1755 -3265
rect 1685 -3295 1695 -3275
rect 1745 -3295 1755 -3275
rect 1685 -3305 1755 -3295
rect 1790 -3275 2020 -3265
rect 1790 -3295 1800 -3275
rect 1830 -3295 1980 -3275
rect 2010 -3295 2020 -3275
rect 1790 -3305 2020 -3295
rect 2485 -3275 2555 -3265
rect 2485 -3295 2495 -3275
rect 2545 -3295 2555 -3275
rect 2485 -3305 2555 -3295
rect 2590 -3275 2820 -3265
rect 2590 -3295 2600 -3275
rect 2630 -3295 2780 -3275
rect 2810 -3295 2820 -3275
rect 2590 -3305 2820 -3295
rect 3285 -3275 3355 -3265
rect 3285 -3295 3295 -3275
rect 3345 -3295 3355 -3275
rect 3285 -3305 3355 -3295
rect 3390 -3275 3620 -3265
rect 3390 -3295 3400 -3275
rect 3430 -3295 3580 -3275
rect 3610 -3295 3620 -3275
rect 3390 -3305 3620 -3295
rect 4085 -3275 4155 -3265
rect 4085 -3295 4095 -3275
rect 4145 -3295 4155 -3275
rect 4085 -3305 4155 -3295
rect 4190 -3275 4420 -3265
rect 4190 -3295 4200 -3275
rect 4230 -3295 4380 -3275
rect 4410 -3295 4420 -3275
rect 4190 -3305 4420 -3295
rect 4885 -3275 4955 -3265
rect 4885 -3295 4895 -3275
rect 4945 -3295 4955 -3275
rect 4885 -3305 4955 -3295
rect 4990 -3275 5220 -3265
rect 4990 -3295 5000 -3275
rect 5030 -3295 5180 -3275
rect 5210 -3295 5220 -3275
rect 4990 -3305 5220 -3295
rect 5790 -3275 5860 -3265
rect 5790 -3295 5800 -3275
rect 5850 -3295 5860 -3275
rect 5790 -3305 5860 -3295
rect 5895 -3270 5945 -3265
rect 6075 -3270 6125 -3265
rect 5895 -3275 6125 -3270
rect 5895 -3295 5905 -3275
rect 5935 -3295 6085 -3275
rect 6115 -3295 6125 -3275
rect 5895 -3305 6125 -3295
rect 6760 -3275 6830 -3265
rect 6760 -3295 6770 -3275
rect 6820 -3295 6830 -3275
rect 6760 -3305 6830 -3295
rect 6690 -4740 6730 -4730
rect 225 -4870 260 -4760
rect 430 -4815 460 -4760
rect 430 -4825 500 -4815
rect 430 -4845 440 -4825
rect 490 -4845 500 -4825
rect 430 -4855 500 -4845
rect 920 -4820 1060 -4790
rect 1230 -4815 1260 -4760
rect 920 -4870 955 -4820
rect 1230 -4825 1300 -4815
rect 1230 -4845 1240 -4825
rect 1290 -4845 1300 -4825
rect 1230 -4855 1300 -4845
rect 1720 -4820 1860 -4790
rect 2030 -4815 2060 -4760
rect 1720 -4870 1755 -4820
rect 2030 -4825 2100 -4815
rect 2030 -4845 2040 -4825
rect 2090 -4845 2100 -4825
rect 2030 -4855 2100 -4845
rect 2520 -4820 2660 -4790
rect 2830 -4815 2860 -4760
rect 2520 -4870 2555 -4820
rect 2830 -4825 2900 -4815
rect 2830 -4845 2840 -4825
rect 2890 -4845 2900 -4825
rect 2830 -4855 2900 -4845
rect 3320 -4820 3460 -4790
rect 3630 -4815 3660 -4760
rect 3320 -4870 3355 -4820
rect 3630 -4825 3700 -4815
rect 3630 -4845 3640 -4825
rect 3690 -4845 3700 -4825
rect 3630 -4855 3700 -4845
rect 4120 -4820 4260 -4790
rect 4430 -4815 4460 -4760
rect 4120 -4870 4155 -4820
rect 4430 -4825 4500 -4815
rect 4430 -4845 4440 -4825
rect 4490 -4845 4500 -4825
rect 4430 -4855 4500 -4845
rect 5025 -4870 5060 -4800
rect 5230 -4815 5260 -4760
rect 5185 -4825 5260 -4815
rect 5185 -4845 5195 -4825
rect 5245 -4845 5260 -4825
rect 5185 -4855 5260 -4845
rect 5825 -4820 5965 -4790
rect 6135 -4815 6165 -4745
rect 6600 -4770 6670 -4760
rect 6600 -4790 6610 -4770
rect 6660 -4790 6670 -4770
rect 6600 -4800 6670 -4790
rect 5825 -4870 5860 -4820
rect 6135 -4825 6205 -4815
rect 6135 -4845 6145 -4825
rect 6195 -4845 6205 -4825
rect 6135 -4855 6205 -4845
rect 225 -4880 295 -4870
rect 225 -4900 235 -4880
rect 285 -4900 295 -4880
rect 225 -4910 295 -4900
rect 885 -4880 955 -4870
rect 885 -4900 895 -4880
rect 945 -4900 955 -4880
rect 885 -4910 955 -4900
rect 990 -4880 1220 -4870
rect 990 -4900 1000 -4880
rect 1030 -4900 1180 -4880
rect 1210 -4900 1220 -4880
rect 990 -4910 1220 -4900
rect 1685 -4880 1755 -4870
rect 1685 -4900 1695 -4880
rect 1745 -4900 1755 -4880
rect 1685 -4910 1755 -4900
rect 1790 -4880 2020 -4870
rect 1790 -4900 1800 -4880
rect 1830 -4900 1980 -4880
rect 2010 -4900 2020 -4880
rect 1790 -4910 2020 -4900
rect 2485 -4880 2555 -4870
rect 2485 -4900 2495 -4880
rect 2545 -4900 2555 -4880
rect 2485 -4910 2555 -4900
rect 2590 -4880 2820 -4870
rect 2590 -4900 2600 -4880
rect 2630 -4900 2780 -4880
rect 2810 -4900 2820 -4880
rect 2590 -4910 2820 -4900
rect 3285 -4880 3355 -4870
rect 3285 -4900 3295 -4880
rect 3345 -4900 3355 -4880
rect 3285 -4910 3355 -4900
rect 3390 -4880 3620 -4870
rect 3390 -4900 3400 -4880
rect 3430 -4900 3580 -4880
rect 3610 -4900 3620 -4880
rect 3390 -4910 3620 -4900
rect 4085 -4880 4155 -4870
rect 4085 -4900 4095 -4880
rect 4145 -4900 4155 -4880
rect 4085 -4910 4155 -4900
rect 4190 -4880 4420 -4870
rect 4190 -4900 4200 -4880
rect 4230 -4900 4380 -4880
rect 4410 -4900 4420 -4880
rect 4190 -4910 4420 -4900
rect 4990 -4880 5060 -4870
rect 4990 -4900 5000 -4880
rect 5050 -4900 5060 -4880
rect 4990 -4910 5060 -4900
rect 5095 -4875 5145 -4870
rect 5275 -4875 5325 -4870
rect 5095 -4880 5325 -4875
rect 5095 -4900 5105 -4880
rect 5135 -4900 5285 -4880
rect 5315 -4900 5325 -4880
rect 5095 -4910 5325 -4900
rect 5790 -4880 5860 -4870
rect 5790 -4900 5800 -4880
rect 5850 -4900 5860 -4880
rect 5790 -4910 5860 -4900
rect 5895 -4880 6125 -4870
rect 5895 -4900 5905 -4880
rect 5935 -4900 6085 -4880
rect 6115 -4900 6125 -4880
rect 5895 -4910 6125 -4900
rect 6630 -4935 6670 -4800
rect 6630 -4985 6640 -4935
rect 6660 -4985 6670 -4935
rect 6630 -4995 6670 -4985
rect 6690 -4790 6700 -4740
rect 6720 -4790 6730 -4740
rect 6690 -4935 6730 -4790
rect 6790 -4740 6830 -4730
rect 6790 -4790 6800 -4740
rect 6820 -4790 6830 -4740
rect 6790 -4870 6830 -4790
rect 6760 -4880 6830 -4870
rect 6760 -4900 6770 -4880
rect 6820 -4900 6830 -4880
rect 6760 -4910 6830 -4900
rect 6690 -4985 6700 -4935
rect 6720 -4985 6730 -4935
rect 6690 -4995 6730 -4985
rect 6630 -6235 6670 -6225
rect 6630 -6285 6640 -6235
rect 6660 -6285 6670 -6235
rect 225 -6475 260 -6365
rect 430 -6420 460 -6365
rect 430 -6430 500 -6420
rect 430 -6450 440 -6430
rect 490 -6450 500 -6430
rect 430 -6460 500 -6450
rect 1025 -6475 1060 -6365
rect 1230 -6420 1260 -6365
rect 1230 -6430 1300 -6420
rect 1230 -6450 1240 -6430
rect 1290 -6450 1300 -6430
rect 1230 -6460 1300 -6450
rect 1825 -6475 1860 -6365
rect 2030 -6420 2060 -6365
rect 2030 -6430 2100 -6420
rect 2030 -6450 2040 -6430
rect 2090 -6450 2100 -6430
rect 2030 -6460 2100 -6450
rect 2625 -6475 2660 -6365
rect 2830 -6420 2860 -6365
rect 2830 -6430 2900 -6420
rect 2830 -6450 2840 -6430
rect 2890 -6450 2900 -6430
rect 2830 -6460 2900 -6450
rect 3425 -6475 3460 -6365
rect 3630 -6420 3660 -6365
rect 3630 -6430 3700 -6420
rect 3630 -6450 3640 -6430
rect 3690 -6450 3700 -6430
rect 3630 -6460 3700 -6450
rect 4225 -6475 4260 -6365
rect 4430 -6420 4460 -6365
rect 4430 -6430 4500 -6420
rect 4430 -6450 4440 -6430
rect 4490 -6450 4500 -6430
rect 4430 -6460 4500 -6450
rect 5130 -6475 5165 -6355
rect 5335 -6420 5365 -6355
rect 5335 -6430 5405 -6420
rect 5335 -6450 5345 -6430
rect 5395 -6450 5405 -6430
rect 5335 -6460 5405 -6450
rect 5930 -6475 5965 -6365
rect 6135 -6420 6165 -6355
rect 6630 -6365 6670 -6285
rect 6600 -6375 6670 -6365
rect 6600 -6395 6610 -6375
rect 6660 -6395 6670 -6375
rect 6600 -6405 6670 -6395
rect 6135 -6430 6205 -6420
rect 6135 -6450 6145 -6430
rect 6195 -6450 6205 -6430
rect 6135 -6460 6205 -6450
rect 225 -6485 295 -6475
rect 225 -6505 235 -6485
rect 285 -6505 295 -6485
rect 225 -6515 295 -6505
rect 1025 -6485 1095 -6475
rect 1025 -6505 1035 -6485
rect 1085 -6505 1095 -6485
rect 1025 -6515 1095 -6505
rect 1825 -6485 1895 -6475
rect 1825 -6505 1835 -6485
rect 1885 -6505 1895 -6485
rect 1825 -6515 1895 -6505
rect 2625 -6485 2695 -6475
rect 2625 -6505 2635 -6485
rect 2685 -6505 2695 -6485
rect 2625 -6515 2695 -6505
rect 3425 -6485 3495 -6475
rect 3425 -6505 3435 -6485
rect 3485 -6505 3495 -6485
rect 3425 -6515 3495 -6505
rect 4225 -6485 4295 -6475
rect 4225 -6505 4235 -6485
rect 4285 -6505 4295 -6485
rect 4225 -6515 4295 -6505
rect 5130 -6485 5200 -6475
rect 5130 -6505 5140 -6485
rect 5190 -6505 5200 -6485
rect 5130 -6515 5200 -6505
rect 5930 -6485 6000 -6475
rect 5930 -6505 5940 -6485
rect 5990 -6505 6000 -6485
rect 5930 -6515 6000 -6505
rect 6630 -6530 6670 -6405
rect 6600 -6540 6670 -6530
rect 6600 -6560 6610 -6540
rect 6660 -6560 6670 -6540
rect 6600 -6570 6670 -6560
rect 6690 -6345 6730 -6335
rect 6690 -6395 6700 -6345
rect 6720 -6395 6730 -6345
rect 6690 -6565 6730 -6395
rect 6790 -6345 6830 -6335
rect 6790 -6395 6800 -6345
rect 6820 -6395 6830 -6345
rect 6790 -6475 6830 -6395
rect 6760 -6485 6830 -6475
rect 6760 -6505 6770 -6485
rect 6820 -6505 6830 -6485
rect 6760 -6515 6830 -6505
rect 6690 -6615 6700 -6565
rect 6720 -6615 6730 -6565
rect 6690 -6625 6730 -6615
<< viali >>
rect 6635 125 6655 175
rect 440 -40 490 -20
rect 1240 -40 1290 -20
rect 2040 -40 2090 -20
rect 2840 -40 2890 -20
rect 3640 -40 3690 -20
rect 4440 -40 4490 -20
rect 5245 -40 5295 -20
rect 6605 20 6655 40
rect 6145 -40 6195 -20
rect 6605 -40 6655 -20
rect 6825 -40 6875 -20
rect 235 -95 285 -75
rect 895 -95 945 -75
rect 1695 -95 1745 -75
rect 2495 -95 2545 -75
rect 3295 -95 3345 -75
rect 4095 -95 4145 -75
rect 4895 -95 4945 -75
rect 5800 -95 5850 -75
rect 6635 -135 6655 -85
rect 6800 -165 6820 -115
rect 6635 -1530 6655 -1480
rect 6745 -1495 6765 -1445
rect 440 -1640 490 -1620
rect 1240 -1640 1290 -1620
rect 2040 -1640 2090 -1620
rect 2840 -1640 2890 -1620
rect 3640 -1640 3690 -1620
rect 4440 -1640 4490 -1620
rect 5240 -1640 5290 -1620
rect 6045 -1640 6095 -1620
rect 6800 -1585 6820 -1535
rect 235 -1695 285 -1675
rect 895 -1695 945 -1675
rect 1695 -1695 1745 -1675
rect 2495 -1695 2545 -1675
rect 3295 -1695 3345 -1675
rect 4095 -1695 4145 -1675
rect 4895 -1695 4945 -1675
rect 5695 -1695 5745 -1675
rect 6770 -1695 6820 -1675
rect 440 -3240 490 -3220
rect 1240 -3240 1290 -3220
rect 2040 -3240 2090 -3220
rect 2840 -3240 2890 -3220
rect 3640 -3240 3690 -3220
rect 4440 -3240 4490 -3220
rect 5240 -3240 5290 -3220
rect 5995 -3240 6045 -3220
rect 6800 -3185 6820 -3135
rect 235 -3295 285 -3275
rect 895 -3295 945 -3275
rect 1695 -3295 1745 -3275
rect 2495 -3295 2545 -3275
rect 3295 -3295 3345 -3275
rect 4095 -3295 4145 -3275
rect 4895 -3295 4945 -3275
rect 5800 -3295 5850 -3275
rect 6770 -3295 6820 -3275
rect 440 -4845 490 -4825
rect 1240 -4845 1290 -4825
rect 2040 -4845 2090 -4825
rect 2840 -4845 2890 -4825
rect 3640 -4845 3690 -4825
rect 4440 -4845 4490 -4825
rect 5195 -4845 5245 -4825
rect 6610 -4790 6660 -4770
rect 6145 -4845 6195 -4825
rect 235 -4900 285 -4880
rect 895 -4900 945 -4880
rect 1695 -4900 1745 -4880
rect 2495 -4900 2545 -4880
rect 3295 -4900 3345 -4880
rect 4095 -4900 4145 -4880
rect 5000 -4900 5050 -4880
rect 5800 -4900 5850 -4880
rect 6640 -4985 6660 -4935
rect 6700 -4790 6720 -4740
rect 6800 -4790 6820 -4740
rect 6770 -4900 6820 -4880
rect 6700 -4985 6720 -4935
rect 6640 -6285 6660 -6235
rect 440 -6450 490 -6430
rect 1240 -6450 1290 -6430
rect 2040 -6450 2090 -6430
rect 2840 -6450 2890 -6430
rect 3640 -6450 3690 -6430
rect 4440 -6450 4490 -6430
rect 5345 -6450 5395 -6430
rect 6610 -6395 6660 -6375
rect 6145 -6450 6195 -6430
rect 235 -6505 285 -6485
rect 1035 -6505 1085 -6485
rect 1835 -6505 1885 -6485
rect 2635 -6505 2685 -6485
rect 3435 -6505 3485 -6485
rect 4235 -6505 4285 -6485
rect 5140 -6505 5190 -6485
rect 5940 -6505 5990 -6485
rect 6610 -6560 6660 -6540
rect 6700 -6395 6720 -6345
rect 6800 -6395 6820 -6345
rect 6770 -6505 6820 -6485
rect 6700 -6615 6720 -6565
<< metal1 >>
rect 0 1545 6775 1585
rect 0 1490 6665 1530
rect 4845 135 4945 1430
rect 6625 175 6665 1490
rect 6625 125 6635 175
rect 6655 125 6665 175
rect 6625 115 6665 125
rect 6735 100 6775 1545
rect 0 60 70 100
rect 6560 60 6775 100
rect 0 5 70 45
rect 6560 40 6720 45
rect 6560 20 6605 40
rect 6655 20 6720 40
rect 6560 5 6720 20
rect 430 -20 6665 -10
rect 430 -40 440 -20
rect 490 -40 1240 -20
rect 1290 -40 2040 -20
rect 2090 -40 2840 -20
rect 2890 -40 3640 -20
rect 3690 -40 4440 -20
rect 4490 -40 5245 -20
rect 5295 -40 6145 -20
rect 6195 -40 6605 -20
rect 6655 -40 6665 -20
rect 430 -50 6665 -40
rect 225 -75 6665 -65
rect 225 -95 235 -75
rect 285 -95 895 -75
rect 945 -95 1695 -75
rect 1745 -95 2495 -75
rect 2545 -95 3295 -75
rect 3345 -95 4095 -75
rect 4145 -95 4895 -75
rect 4945 -95 5800 -75
rect 5850 -85 6665 -75
rect 5850 -95 6635 -85
rect 225 -105 6635 -95
rect 6625 -135 6635 -105
rect 6655 -135 6665 -85
rect 6625 -145 6665 -135
rect 5635 -1465 5755 -170
rect 6625 -1480 6665 -1470
rect 6625 -1500 6635 -1480
rect 0 -1540 70 -1500
rect 6555 -1530 6635 -1500
rect 6655 -1530 6665 -1480
rect 6555 -1540 6665 -1530
rect 6680 -1555 6720 5
rect 6735 -1445 6775 60
rect 6815 -20 6885 -10
rect 6815 -40 6825 -20
rect 6875 -40 6885 -20
rect 6815 -50 6885 -40
rect 6735 -1495 6745 -1445
rect 6765 -1495 6775 -1445
rect 6735 -1505 6775 -1495
rect 6790 -115 6830 -105
rect 6790 -165 6800 -115
rect 6820 -165 6830 -115
rect 0 -1595 70 -1555
rect 6555 -1595 6720 -1555
rect 6790 -1535 6830 -165
rect 6790 -1585 6800 -1535
rect 6820 -1585 6830 -1535
rect 6790 -1595 6830 -1585
rect 6845 -1610 6885 -50
rect 430 -1620 6885 -1610
rect 430 -1640 440 -1620
rect 490 -1640 1240 -1620
rect 1290 -1640 2040 -1620
rect 2090 -1640 2840 -1620
rect 2890 -1640 3640 -1620
rect 3690 -1640 4440 -1620
rect 4490 -1640 5240 -1620
rect 5290 -1640 6045 -1620
rect 6095 -1640 6885 -1620
rect 430 -1650 6885 -1640
rect 225 -1675 6830 -1665
rect 225 -1695 235 -1675
rect 285 -1695 895 -1675
rect 945 -1695 1695 -1675
rect 1745 -1695 2495 -1675
rect 2545 -1695 3295 -1675
rect 3345 -1695 4095 -1675
rect 4145 -1695 4895 -1675
rect 4945 -1695 5695 -1675
rect 5745 -1695 6770 -1675
rect 6820 -1695 6830 -1675
rect 225 -1705 6830 -1695
rect 0 -3140 70 -3100
rect 6790 -3135 6830 -1705
rect 0 -3195 70 -3155
rect 6790 -3185 6800 -3135
rect 6820 -3185 6830 -3135
rect 6790 -3195 6830 -3185
rect 6845 -3210 6885 -1650
rect 430 -3220 6885 -3210
rect 430 -3240 440 -3220
rect 490 -3240 1240 -3220
rect 1290 -3240 2040 -3220
rect 2090 -3240 2840 -3220
rect 2890 -3240 3640 -3220
rect 3690 -3240 4440 -3220
rect 4490 -3240 5240 -3220
rect 5290 -3240 5995 -3220
rect 6045 -3240 6885 -3220
rect 430 -3250 6885 -3240
rect 225 -3275 6830 -3265
rect 225 -3295 235 -3275
rect 285 -3295 895 -3275
rect 945 -3295 1695 -3275
rect 1745 -3295 2495 -3275
rect 2545 -3295 3295 -3275
rect 3345 -3295 4095 -3275
rect 4145 -3295 4895 -3275
rect 4945 -3295 5800 -3275
rect 5850 -3295 6770 -3275
rect 6820 -3295 6830 -3275
rect 225 -3305 6830 -3295
rect 5635 -4670 5765 -3375
rect 0 -4745 70 -4705
rect 6565 -4740 6730 -4705
rect 6565 -4745 6700 -4740
rect 0 -4800 70 -4760
rect 6565 -4770 6670 -4760
rect 6565 -4790 6610 -4770
rect 6660 -4790 6670 -4770
rect 6565 -4800 6670 -4790
rect 6690 -4790 6700 -4745
rect 6720 -4790 6730 -4740
rect 6690 -4800 6730 -4790
rect 6790 -4740 6830 -3305
rect 6790 -4790 6800 -4740
rect 6820 -4790 6830 -4740
rect 6790 -4800 6830 -4790
rect 6845 -4815 6885 -3250
rect 430 -4825 6885 -4815
rect 430 -4845 440 -4825
rect 490 -4845 1240 -4825
rect 1290 -4845 2040 -4825
rect 2090 -4845 2840 -4825
rect 2890 -4845 3640 -4825
rect 3690 -4845 4440 -4825
rect 4490 -4845 5195 -4825
rect 5245 -4845 6145 -4825
rect 6195 -4845 6885 -4825
rect 430 -4855 6885 -4845
rect 225 -4880 6830 -4870
rect 225 -4900 235 -4880
rect 285 -4900 895 -4880
rect 945 -4900 1695 -4880
rect 1745 -4900 2495 -4880
rect 2545 -4900 3295 -4880
rect 3345 -4900 4095 -4880
rect 4145 -4900 5000 -4880
rect 5050 -4900 5800 -4880
rect 5850 -4900 6770 -4880
rect 6820 -4900 6830 -4880
rect 225 -4910 6830 -4900
rect 6630 -4935 6670 -4925
rect 4835 -6275 4950 -4980
rect 6630 -4985 6640 -4935
rect 6660 -4985 6670 -4935
rect 6630 -6235 6670 -4985
rect 6630 -6285 6640 -6235
rect 6660 -6285 6670 -6235
rect 6630 -6295 6670 -6285
rect 6690 -4935 6730 -4925
rect 6690 -4985 6700 -4935
rect 6720 -4985 6730 -4935
rect 6690 -6310 6730 -4985
rect 0 -6350 70 -6310
rect 6560 -6345 6730 -6310
rect 6560 -6350 6700 -6345
rect 0 -6405 70 -6365
rect 6560 -6375 6670 -6365
rect 6560 -6395 6610 -6375
rect 6660 -6395 6670 -6375
rect 6560 -6405 6670 -6395
rect 6690 -6395 6700 -6350
rect 6720 -6395 6730 -6345
rect 6690 -6405 6730 -6395
rect 6790 -6345 6830 -4910
rect 6790 -6395 6800 -6345
rect 6820 -6395 6830 -6345
rect 6790 -6405 6830 -6395
rect 6845 -6420 6885 -4855
rect 430 -6430 6885 -6420
rect 430 -6450 440 -6430
rect 490 -6450 1240 -6430
rect 1290 -6450 2040 -6430
rect 2090 -6450 2840 -6430
rect 2890 -6450 3640 -6430
rect 3690 -6450 4440 -6430
rect 4490 -6450 5345 -6430
rect 5395 -6450 6145 -6430
rect 6195 -6450 6885 -6430
rect 430 -6460 6885 -6450
rect 225 -6485 6830 -6475
rect 225 -6505 235 -6485
rect 285 -6505 1035 -6485
rect 1085 -6505 1835 -6485
rect 1885 -6505 2635 -6485
rect 2685 -6505 3435 -6485
rect 3485 -6505 4235 -6485
rect 4285 -6505 5140 -6485
rect 5190 -6505 5940 -6485
rect 5990 -6505 6770 -6485
rect 6820 -6505 6830 -6485
rect 225 -6515 6830 -6505
rect 0 -6540 6670 -6530
rect 0 -6560 6610 -6540
rect 6660 -6560 6670 -6540
rect 0 -6570 6670 -6560
rect 6690 -6565 6730 -6555
rect 6690 -6585 6700 -6565
rect 0 -6615 6700 -6585
rect 6720 -6615 6730 -6565
rect 0 -6625 6730 -6615
rect 6790 -6585 6830 -6515
rect 6845 -6505 6885 -6460
rect 6845 -6545 6890 -6505
rect 6790 -6625 6890 -6585
use dac_unit  dac_unit_0
timestamp 1702614989
transform 1 0 -1115 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_1
timestamp 1702614989
transform 1 0 -315 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_2
timestamp 1702614989
transform 1 0 485 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_3
timestamp 1702614989
transform 1 0 1285 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_4
timestamp 1702614989
transform 1 0 2085 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_5
timestamp 1702614989
transform 1 0 4590 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_6
timestamp 1702614989
transform 1 0 -1115 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_7
timestamp 1702614989
transform 1 0 2085 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_8
timestamp 1702614989
transform 1 0 -315 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_9
timestamp 1702614989
transform 1 0 485 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_10
timestamp 1702614989
transform 1 0 1285 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_11
timestamp 1702614989
transform 1 0 4485 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_12
timestamp 1702614989
transform 1 0 2885 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_13
timestamp 1702614989
transform 1 0 -1115 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_14
timestamp 1702614989
transform 1 0 3685 0 1 -3250
box 1115 55 2005 1520
use dac_unit  dac_unit_15
timestamp 1702614989
transform 1 0 -315 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_16
timestamp 1702614989
transform 1 0 485 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_17
timestamp 1702614989
transform 1 0 1285 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_18
timestamp 1702614989
transform 1 0 2085 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_19
timestamp 1702614989
transform 1 0 2885 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_20
timestamp 1702614989
transform 1 0 3685 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_21
timestamp 1702614989
transform 1 0 -1115 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_22
timestamp 1702614989
transform 1 0 -315 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_23
timestamp 1702614989
transform 1 0 485 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_24
timestamp 1702614989
transform 1 0 1285 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_25
timestamp 1702614989
transform 1 0 2885 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_26
timestamp 1702614989
transform 1 0 -1115 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_27
timestamp 1702614989
transform 1 0 3685 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_28
timestamp 1702614989
transform 1 0 2085 0 1 -1650
box 1115 55 2005 1520
use dac_unit  dac_unit_29
timestamp 1702614989
transform 1 0 2885 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_30
timestamp 1702614989
transform 1 0 2885 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_31
timestamp 1702614989
transform 1 0 2085 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_32
timestamp 1702614989
transform 1 0 1285 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_33
timestamp 1702614989
transform 1 0 485 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_34
timestamp 1702614989
transform 1 0 -315 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_35
timestamp 1702614989
transform 1 0 3790 0 1 -50
box 1115 55 2005 1520
use dac_unit  dac_unit_36
timestamp 1702614989
transform 1 0 3790 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_37
timestamp 1702614989
transform 1 0 4590 0 1 -6460
box 1115 55 2005 1520
use dac_unit  dac_unit_38
timestamp 1702614989
transform 1 0 4590 0 1 -4855
box 1115 55 2005 1520
use dac_unit  dac_unit_40
timestamp 1702614989
transform 1 0 4590 0 1 -50
box 1115 55 2005 1520
<< labels >>
rlabel metal1 6890 -6525 6890 -6525 3 Viout-
rlabel metal1 6890 -6605 6890 -6605 3 Viout+
rlabel metal1 0 1560 0 1560 7 Vphi1
rlabel metal1 0 1510 0 1510 7 Vphi1_b
rlabel metal1 0 80 0 80 7 Vphi2
rlabel metal1 0 25 0 25 7 Vphi2_b
rlabel metal1 0 -1520 0 -1520 7 Vphi3
rlabel metal1 0 -1575 0 -1575 7 Vphi3_b
rlabel metal1 0 -3120 0 -3120 7 Vphi4
rlabel metal1 0 -3175 0 -3175 7 Vphi4_b
rlabel metal1 0 -4725 0 -4725 7 Vphi5
rlabel metal1 0 -4780 0 -4780 7 Vphi5_b
rlabel metal1 0 -6330 0 -6330 7 Vphi6
rlabel metal1 0 -6385 0 -6385 7 Vphi6_b
rlabel poly 6000 1585 6000 1585 1 Vbp
rlabel poly 6100 1585 6100 1585 1 Vcp
rlabel metal1 0 -6550 0 -6550 7 Vphi7_b
rlabel metal1 0 -6605 0 -6605 7 Vphi7
<< end >>
