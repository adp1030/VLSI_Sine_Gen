magic
tech sky130A
timestamp 1702516191
<< nwell >>
rect 6420 -145 6460 -90
rect 6335 -175 6460 -145
rect -30 -315 0 -175
rect 6420 -230 6460 -175
rect 6670 -230 6700 -90
rect -30 -2240 0 -2100
rect -30 -4165 0 -4025
rect -30 -6090 0 -5950
rect -30 -8015 0 -7875
rect 6420 -8015 6460 -7875
rect 6670 -8015 6700 -7875
<< poly >>
rect -340 15 9080 25
rect -340 -5 -330 15
rect -310 10 9080 15
rect -310 -5 -300 10
rect -340 -15 -300 -5
rect -380 -50 -340 -40
rect -380 -70 -370 -50
rect -350 -65 -340 -50
rect -240 -50 -200 -40
rect -240 -65 -230 -50
rect -350 -70 -230 -65
rect -210 -70 -200 -50
rect -380 -80 -200 -70
rect 6925 -55 6940 10
rect 7995 -55 8010 10
rect 9065 -55 9080 10
rect 6925 -65 6975 -55
rect 6925 -85 6935 -65
rect 6955 -85 6975 -65
rect 6925 -90 6975 -85
rect 7995 -65 8045 -55
rect 7995 -85 8005 -65
rect 8025 -85 8045 -65
rect 7995 -90 8045 -85
rect 9065 -65 9115 -55
rect 9065 -85 9075 -65
rect 9095 -85 9115 -65
rect 9065 -90 9115 -85
rect -340 -150 275 -140
rect -340 -170 -330 -150
rect -310 -155 235 -150
rect -310 -170 -300 -155
rect -340 -180 -300 -170
rect 225 -170 235 -155
rect 255 -160 275 -150
rect 1295 -150 1345 -140
rect 1295 -160 1305 -150
rect 255 -170 1305 -160
rect 1325 -160 1345 -150
rect 2365 -150 2415 -140
rect 2365 -160 2375 -150
rect 1325 -170 2375 -160
rect 2395 -160 2415 -150
rect 3435 -150 3485 -140
rect 3435 -160 3445 -150
rect 2395 -170 3445 -160
rect 3465 -160 3485 -150
rect 4505 -150 4555 -140
rect 4505 -160 4515 -150
rect 3465 -170 4515 -160
rect 4535 -160 4555 -150
rect 5575 -150 5625 -140
rect 5575 -160 5585 -150
rect 4535 -170 5585 -160
rect 5605 -170 5625 -150
rect 225 -175 5625 -170
rect -380 -1160 -340 -1150
rect -380 -1180 -370 -1160
rect -350 -1175 -340 -1160
rect -240 -1160 -200 -1150
rect -240 -1175 -230 -1160
rect -350 -1180 -230 -1175
rect -210 -1180 -200 -1160
rect -380 -1190 -200 -1180
rect 7125 -1850 7165 -1840
rect 7125 -1870 7135 -1850
rect 7155 -1865 7165 -1850
rect 8195 -1850 8235 -1840
rect 8195 -1865 8205 -1850
rect 7155 -1870 8205 -1865
rect 8225 -1865 8235 -1850
rect 9265 -1850 9305 -1840
rect 9265 -1865 9275 -1850
rect 8225 -1870 9275 -1865
rect 9295 -1865 9305 -1850
rect 9295 -1870 9925 -1865
rect 7125 -1880 9925 -1870
rect 425 -1935 465 -1925
rect 425 -1955 435 -1935
rect 455 -1950 465 -1935
rect 1495 -1935 1535 -1925
rect 1495 -1950 1505 -1935
rect 455 -1955 1505 -1950
rect 1525 -1950 1535 -1935
rect 2565 -1935 2605 -1925
rect 2565 -1950 2575 -1935
rect 1525 -1955 2575 -1950
rect 2595 -1950 2605 -1935
rect 3635 -1935 3675 -1925
rect 3635 -1950 3645 -1935
rect 2595 -1955 3645 -1950
rect 3665 -1950 3675 -1935
rect 4705 -1935 4745 -1925
rect 4705 -1950 4715 -1935
rect 3665 -1955 4715 -1950
rect 4735 -1950 4745 -1935
rect 5775 -1935 5815 -1925
rect 5775 -1950 5785 -1935
rect 4735 -1955 5785 -1950
rect 5805 -1950 5815 -1935
rect 9910 -1950 9925 -1880
rect 5805 -1955 9925 -1950
rect 425 -1965 9925 -1955
rect -340 -2075 275 -2065
rect -340 -2095 -330 -2075
rect -310 -2080 235 -2075
rect -310 -2095 -300 -2080
rect -340 -2105 -300 -2095
rect 225 -2095 235 -2080
rect 255 -2085 275 -2075
rect 1295 -2075 1345 -2065
rect 1295 -2085 1305 -2075
rect 255 -2095 1305 -2085
rect 1325 -2085 1345 -2075
rect 2365 -2075 2415 -2065
rect 2365 -2085 2375 -2075
rect 1325 -2095 2375 -2085
rect 2395 -2085 2415 -2075
rect 3435 -2075 3485 -2065
rect 3435 -2085 3445 -2075
rect 2395 -2095 3445 -2085
rect 3465 -2085 3485 -2075
rect 4505 -2075 4555 -2065
rect 4505 -2085 4515 -2075
rect 3465 -2095 4515 -2085
rect 4535 -2085 4555 -2075
rect 5575 -2075 5625 -2065
rect 5575 -2085 5585 -2075
rect 4535 -2095 5585 -2085
rect 5605 -2085 5625 -2075
rect 6645 -2075 6695 -2065
rect 6645 -2085 6655 -2075
rect 5605 -2095 6655 -2085
rect 6675 -2085 6695 -2075
rect 6675 -2095 7490 -2085
rect 225 -2100 7490 -2095
rect -380 -3085 -340 -3075
rect -380 -3105 -370 -3085
rect -350 -3100 -340 -3085
rect -240 -3085 -200 -3075
rect -240 -3100 -230 -3085
rect -350 -3105 -230 -3100
rect -210 -3105 -200 -3085
rect -380 -3115 -200 -3105
rect 425 -3860 465 -3850
rect 425 -3880 435 -3860
rect 455 -3875 465 -3860
rect 1495 -3860 1535 -3850
rect 1495 -3875 1505 -3860
rect 455 -3880 1505 -3875
rect 1525 -3875 1535 -3860
rect 2565 -3860 2605 -3850
rect 2565 -3875 2575 -3860
rect 1525 -3880 2575 -3875
rect 2595 -3875 2605 -3860
rect 3635 -3860 3675 -3850
rect 3635 -3875 3645 -3860
rect 2595 -3880 3645 -3875
rect 3665 -3875 3675 -3860
rect 4705 -3860 4745 -3850
rect 4705 -3875 4715 -3860
rect 3665 -3880 4715 -3875
rect 4735 -3875 4745 -3860
rect 5775 -3860 5815 -3850
rect 5775 -3875 5785 -3860
rect 4735 -3880 5785 -3875
rect 5805 -3875 5815 -3860
rect 6845 -3860 6885 -3850
rect 6845 -3875 6855 -3860
rect 5805 -3880 6855 -3875
rect 6875 -3875 6885 -3860
rect 9910 -3875 9925 -1965
rect 6875 -3880 9925 -3875
rect 425 -3890 9925 -3880
rect -340 -4000 275 -3990
rect -340 -4020 -330 -4000
rect -310 -4005 235 -4000
rect -310 -4020 -300 -4005
rect -340 -4030 -300 -4020
rect 225 -4020 235 -4005
rect 255 -4010 275 -4000
rect 1295 -4000 1345 -3990
rect 1295 -4010 1305 -4000
rect 255 -4020 1305 -4010
rect 1325 -4010 1345 -4000
rect 2365 -4000 2415 -3990
rect 2365 -4010 2375 -4000
rect 1325 -4020 2375 -4010
rect 2395 -4010 2415 -4000
rect 3435 -4000 3485 -3990
rect 3435 -4010 3445 -4000
rect 2395 -4020 3445 -4010
rect 3465 -4010 3485 -4000
rect 4505 -4000 4555 -3990
rect 4505 -4010 4515 -4000
rect 3465 -4020 4515 -4010
rect 4535 -4010 4555 -4000
rect 5575 -4000 5625 -3990
rect 5575 -4010 5585 -4000
rect 4535 -4020 5585 -4010
rect 5605 -4010 5625 -4000
rect 6645 -4000 6695 -3990
rect 6645 -4010 6655 -4000
rect 5605 -4020 6655 -4010
rect 6675 -4010 6695 -4000
rect 7715 -4000 7765 -3990
rect 7715 -4010 7725 -4000
rect 6675 -4020 7725 -4010
rect 7745 -4020 7765 -4000
rect 225 -4025 7765 -4020
rect -380 -5010 -340 -5000
rect -380 -5030 -370 -5010
rect -350 -5025 -340 -5010
rect -240 -5010 -200 -5000
rect -240 -5025 -230 -5010
rect -350 -5030 -230 -5025
rect -210 -5030 -200 -5010
rect -380 -5040 -200 -5030
rect 425 -5785 465 -5775
rect 425 -5805 435 -5785
rect 455 -5800 465 -5785
rect 1495 -5785 1535 -5775
rect 1495 -5800 1505 -5785
rect 455 -5805 1505 -5800
rect 1525 -5800 1535 -5785
rect 2565 -5785 2605 -5775
rect 2565 -5800 2575 -5785
rect 1525 -5805 2575 -5800
rect 2595 -5800 2605 -5785
rect 3635 -5785 3675 -5775
rect 3635 -5800 3645 -5785
rect 2595 -5805 3645 -5800
rect 3665 -5800 3675 -5785
rect 4705 -5785 4745 -5775
rect 4705 -5800 4715 -5785
rect 3665 -5805 4715 -5800
rect 4735 -5800 4745 -5785
rect 5775 -5785 5815 -5775
rect 5775 -5800 5785 -5785
rect 4735 -5805 5785 -5800
rect 5805 -5800 5815 -5785
rect 6845 -5785 6885 -5775
rect 6845 -5800 6855 -5785
rect 5805 -5805 6855 -5800
rect 6875 -5800 6885 -5785
rect 7915 -5785 7955 -5775
rect 7915 -5800 7925 -5785
rect 6875 -5805 7925 -5800
rect 7945 -5800 7955 -5785
rect 9910 -5800 9925 -3890
rect 7945 -5805 9925 -5800
rect 425 -5815 9925 -5805
rect -340 -5925 275 -5915
rect -340 -5945 -330 -5925
rect -310 -5930 235 -5925
rect -310 -5945 -300 -5930
rect -340 -5955 -300 -5945
rect 225 -5945 235 -5930
rect 255 -5935 275 -5925
rect 1295 -5925 1345 -5915
rect 1295 -5935 1305 -5925
rect 255 -5945 1305 -5935
rect 1325 -5935 1345 -5925
rect 2365 -5925 2415 -5915
rect 2365 -5935 2375 -5925
rect 1325 -5945 2375 -5935
rect 2395 -5935 2415 -5925
rect 3435 -5925 3485 -5915
rect 3435 -5935 3445 -5925
rect 2395 -5945 3445 -5935
rect 3465 -5935 3485 -5925
rect 4505 -5925 4555 -5915
rect 4505 -5935 4515 -5925
rect 3465 -5945 4515 -5935
rect 4535 -5935 4555 -5925
rect 5575 -5925 5625 -5915
rect 5575 -5935 5585 -5925
rect 4535 -5945 5585 -5935
rect 5605 -5935 5625 -5925
rect 6645 -5925 6695 -5915
rect 6645 -5935 6655 -5925
rect 5605 -5945 6655 -5935
rect 6675 -5935 6695 -5925
rect 6675 -5945 7490 -5935
rect 225 -5950 7490 -5945
rect -380 -6935 -340 -6925
rect -380 -6955 -370 -6935
rect -350 -6950 -340 -6935
rect -240 -6935 -200 -6925
rect -240 -6950 -230 -6935
rect -350 -6955 -230 -6950
rect -210 -6955 -200 -6935
rect -380 -6965 -200 -6955
rect 425 -7710 465 -7700
rect 425 -7730 435 -7710
rect 455 -7725 465 -7710
rect 1495 -7710 1535 -7700
rect 1495 -7725 1505 -7710
rect 455 -7730 1505 -7725
rect 1525 -7725 1535 -7710
rect 2565 -7710 2605 -7700
rect 2565 -7725 2575 -7710
rect 1525 -7730 2575 -7725
rect 2595 -7725 2605 -7710
rect 3635 -7710 3675 -7700
rect 3635 -7725 3645 -7710
rect 2595 -7730 3645 -7725
rect 3665 -7725 3675 -7710
rect 4705 -7710 4745 -7700
rect 4705 -7725 4715 -7710
rect 3665 -7730 4715 -7725
rect 4735 -7725 4745 -7710
rect 5775 -7710 5815 -7700
rect 5775 -7725 5785 -7710
rect 4735 -7730 5785 -7725
rect 5805 -7725 5815 -7710
rect 6845 -7710 6885 -7700
rect 6845 -7725 6855 -7710
rect 5805 -7730 6855 -7725
rect 6875 -7725 6885 -7710
rect 9910 -7725 9925 -5815
rect 6875 -7730 9925 -7725
rect 425 -7740 9925 -7730
rect -340 -7850 275 -7840
rect -340 -7870 -330 -7850
rect -310 -7855 235 -7850
rect -310 -7870 -300 -7855
rect -340 -7880 -300 -7870
rect 225 -7870 235 -7855
rect 255 -7860 275 -7850
rect 1295 -7850 1345 -7840
rect 1295 -7860 1305 -7850
rect 255 -7870 1305 -7860
rect 1325 -7860 1345 -7850
rect 2365 -7850 2415 -7840
rect 2365 -7860 2375 -7850
rect 1325 -7870 2375 -7860
rect 2395 -7860 2415 -7850
rect 3435 -7850 3485 -7840
rect 3435 -7860 3445 -7850
rect 2395 -7870 3445 -7860
rect 3465 -7860 3485 -7850
rect 4505 -7850 4555 -7840
rect 4505 -7860 4515 -7850
rect 3465 -7870 4515 -7860
rect 4535 -7860 4555 -7850
rect 5575 -7850 5625 -7840
rect 5575 -7860 5585 -7850
rect 4535 -7870 5585 -7860
rect 5605 -7860 5625 -7850
rect 6525 -7850 6655 -7835
rect 6525 -7860 6540 -7850
rect 5605 -7870 6540 -7860
rect 225 -7875 6540 -7870
rect 6640 -7860 6655 -7850
rect 6925 -7850 6975 -7840
rect 6925 -7860 6935 -7850
rect 6640 -7870 6935 -7860
rect 6955 -7860 6975 -7850
rect 7995 -7850 8045 -7840
rect 7995 -7860 8005 -7850
rect 6955 -7870 8005 -7860
rect 8025 -7860 8045 -7850
rect 9065 -7850 9115 -7840
rect 9065 -7860 9075 -7850
rect 8025 -7870 9075 -7860
rect 9095 -7870 9115 -7850
rect 6640 -7875 9115 -7870
rect -380 -8860 -340 -8850
rect -380 -8880 -370 -8860
rect -350 -8875 -340 -8860
rect -240 -8860 -200 -8850
rect -240 -8875 -230 -8860
rect -350 -8880 -230 -8875
rect -210 -8880 -200 -8860
rect -380 -8890 -200 -8880
rect 7125 -9635 7165 -9625
rect 7125 -9655 7135 -9635
rect 7155 -9650 7165 -9635
rect 8195 -9635 8235 -9625
rect 8195 -9650 8205 -9635
rect 7155 -9655 8205 -9650
rect 8225 -9650 8235 -9635
rect 9265 -9635 9305 -9625
rect 9265 -9650 9275 -9635
rect 8225 -9655 9275 -9650
rect 9295 -9650 9305 -9635
rect 9910 -9650 9925 -7740
rect 9295 -9655 9925 -9650
rect 7125 -9665 9925 -9655
rect 425 -9710 465 -9700
rect 425 -9730 435 -9710
rect 455 -9725 465 -9710
rect 1495 -9710 1535 -9700
rect 1495 -9725 1505 -9710
rect 455 -9730 1505 -9725
rect 1525 -9725 1535 -9710
rect 2565 -9710 2605 -9700
rect 2565 -9725 2575 -9710
rect 1525 -9730 2575 -9725
rect 2595 -9725 2605 -9710
rect 3635 -9710 3675 -9700
rect 3635 -9725 3645 -9710
rect 2595 -9730 3645 -9725
rect 3665 -9725 3675 -9710
rect 4705 -9710 4745 -9700
rect 4705 -9725 4715 -9710
rect 3665 -9730 4715 -9725
rect 4735 -9725 4745 -9710
rect 5775 -9710 5815 -9700
rect 5775 -9725 5785 -9710
rect 4735 -9730 5785 -9725
rect 5805 -9725 5815 -9710
rect 9910 -9725 9925 -9665
rect 5805 -9730 9925 -9725
rect 425 -9740 9925 -9730
rect 6390 -9775 6735 -9765
rect 6390 -9795 6400 -9775
rect 6420 -9780 6705 -9775
rect 6420 -9795 6430 -9780
rect 6390 -9805 6430 -9795
rect 6695 -9795 6705 -9780
rect 6725 -9795 6735 -9775
rect 6695 -9805 6735 -9795
rect -380 -9815 -340 -9805
rect -380 -9835 -370 -9815
rect -350 -9830 -340 -9815
rect -240 -9815 -200 -9805
rect -240 -9830 -230 -9815
rect -350 -9835 -230 -9830
rect -210 -9835 -200 -9815
rect 9910 -9810 9925 -9740
rect 9985 -9795 10025 -9785
rect 9985 -9810 9995 -9795
rect 9910 -9815 9995 -9810
rect 10015 -9815 10025 -9795
rect 9910 -9825 10025 -9815
rect -380 -9845 -200 -9835
<< polycont >>
rect -330 -5 -310 15
rect -370 -70 -350 -50
rect -230 -70 -210 -50
rect 6935 -85 6955 -65
rect 8005 -85 8025 -65
rect 9075 -85 9095 -65
rect -330 -170 -310 -150
rect 235 -170 255 -150
rect 1305 -170 1325 -150
rect 2375 -170 2395 -150
rect 3445 -170 3465 -150
rect 4515 -170 4535 -150
rect 5585 -170 5605 -150
rect -370 -1180 -350 -1160
rect -230 -1180 -210 -1160
rect 7135 -1870 7155 -1850
rect 8205 -1870 8225 -1850
rect 9275 -1870 9295 -1850
rect 435 -1955 455 -1935
rect 1505 -1955 1525 -1935
rect 2575 -1955 2595 -1935
rect 3645 -1955 3665 -1935
rect 4715 -1955 4735 -1935
rect 5785 -1955 5805 -1935
rect -330 -2095 -310 -2075
rect 235 -2095 255 -2075
rect 1305 -2095 1325 -2075
rect 2375 -2095 2395 -2075
rect 3445 -2095 3465 -2075
rect 4515 -2095 4535 -2075
rect 5585 -2095 5605 -2075
rect 6655 -2095 6675 -2075
rect -370 -3105 -350 -3085
rect -230 -3105 -210 -3085
rect 435 -3880 455 -3860
rect 1505 -3880 1525 -3860
rect 2575 -3880 2595 -3860
rect 3645 -3880 3665 -3860
rect 4715 -3880 4735 -3860
rect 5785 -3880 5805 -3860
rect 6855 -3880 6875 -3860
rect -330 -4020 -310 -4000
rect 235 -4020 255 -4000
rect 1305 -4020 1325 -4000
rect 2375 -4020 2395 -4000
rect 3445 -4020 3465 -4000
rect 4515 -4020 4535 -4000
rect 5585 -4020 5605 -4000
rect 6655 -4020 6675 -4000
rect 7725 -4020 7745 -4000
rect -370 -5030 -350 -5010
rect -230 -5030 -210 -5010
rect 435 -5805 455 -5785
rect 1505 -5805 1525 -5785
rect 2575 -5805 2595 -5785
rect 3645 -5805 3665 -5785
rect 4715 -5805 4735 -5785
rect 5785 -5805 5805 -5785
rect 6855 -5805 6875 -5785
rect 7925 -5805 7945 -5785
rect -330 -5945 -310 -5925
rect 235 -5945 255 -5925
rect 1305 -5945 1325 -5925
rect 2375 -5945 2395 -5925
rect 3445 -5945 3465 -5925
rect 4515 -5945 4535 -5925
rect 5585 -5945 5605 -5925
rect 6655 -5945 6675 -5925
rect -370 -6955 -350 -6935
rect -230 -6955 -210 -6935
rect 435 -7730 455 -7710
rect 1505 -7730 1525 -7710
rect 2575 -7730 2595 -7710
rect 3645 -7730 3665 -7710
rect 4715 -7730 4735 -7710
rect 5785 -7730 5805 -7710
rect 6855 -7730 6875 -7710
rect -330 -7870 -310 -7850
rect 235 -7870 255 -7850
rect 1305 -7870 1325 -7850
rect 2375 -7870 2395 -7850
rect 3445 -7870 3465 -7850
rect 4515 -7870 4535 -7850
rect 5585 -7870 5605 -7850
rect 6935 -7870 6955 -7850
rect 8005 -7870 8025 -7850
rect 9075 -7870 9095 -7850
rect -370 -8880 -350 -8860
rect -230 -8880 -210 -8860
rect 7135 -9655 7155 -9635
rect 8205 -9655 8225 -9635
rect 9275 -9655 9295 -9635
rect 435 -9730 455 -9710
rect 1505 -9730 1525 -9710
rect 2575 -9730 2595 -9710
rect 3645 -9730 3665 -9710
rect 4715 -9730 4735 -9710
rect 5785 -9730 5805 -9710
rect 6400 -9795 6420 -9775
rect 6705 -9795 6725 -9775
rect -370 -9835 -350 -9815
rect -230 -9835 -210 -9815
rect 9995 -9815 10015 -9795
<< locali >>
rect -400 45 9190 65
rect -400 15 -300 25
rect -400 5 -330 15
rect -340 -5 -330 5
rect -310 -5 -300 15
rect -340 -15 -300 -5
rect -380 -50 -340 -40
rect -380 -60 -370 -50
rect -400 -70 -370 -60
rect -350 -70 -340 -50
rect -400 -80 -340 -70
rect -320 -140 -300 -15
rect -340 -150 -300 -140
rect -340 -170 -330 -150
rect -310 -170 -300 -150
rect -340 -180 -300 -170
rect -380 -1160 -340 -1150
rect -380 -1170 -370 -1160
rect -400 -1180 -370 -1170
rect -350 -1180 -340 -1160
rect -400 -1190 -340 -1180
rect -320 -2065 -300 -180
rect -340 -2075 -300 -2065
rect -340 -2095 -330 -2075
rect -310 -2095 -300 -2075
rect -340 -2105 -300 -2095
rect -380 -3085 -340 -3075
rect -380 -3095 -370 -3085
rect -400 -3105 -370 -3095
rect -350 -3105 -340 -3085
rect -400 -3115 -340 -3105
rect -320 -3990 -300 -2105
rect -340 -4000 -300 -3990
rect -340 -4020 -330 -4000
rect -310 -4020 -300 -4000
rect -340 -4030 -300 -4020
rect -380 -5010 -340 -5000
rect -380 -5020 -370 -5010
rect -400 -5030 -370 -5020
rect -350 -5030 -340 -5010
rect -400 -5040 -340 -5030
rect -320 -5915 -300 -4030
rect -340 -5925 -300 -5915
rect -340 -5945 -330 -5925
rect -310 -5945 -300 -5925
rect -340 -5955 -300 -5945
rect -380 -6935 -340 -6925
rect -380 -6945 -370 -6935
rect -400 -6955 -370 -6945
rect -350 -6955 -340 -6935
rect -400 -6965 -340 -6955
rect -320 -7840 -300 -5955
rect -280 -100 -260 45
rect -240 -50 -200 -40
rect -240 -70 -230 -50
rect -210 -60 -200 -50
rect -210 -70 6460 -60
rect -240 -80 6460 -70
rect -280 -120 5700 -100
rect -280 -2025 -260 -120
rect 225 -150 275 -140
rect 225 -170 235 -150
rect 255 -170 275 -150
rect 225 -175 275 -170
rect 330 -175 350 -120
rect 1295 -150 1345 -140
rect 1295 -170 1305 -150
rect 1325 -170 1345 -150
rect 1295 -175 1345 -170
rect 1400 -175 1420 -120
rect 2365 -150 2415 -140
rect 2365 -170 2375 -150
rect 2395 -170 2415 -150
rect 2365 -175 2415 -170
rect 2470 -175 2490 -120
rect 3435 -150 3485 -140
rect 3435 -170 3445 -150
rect 3465 -170 3485 -150
rect 3435 -175 3485 -170
rect 3540 -175 3560 -120
rect 4505 -150 4555 -140
rect 4505 -170 4515 -150
rect 4535 -170 4555 -150
rect 4505 -175 4555 -170
rect 4610 -175 4630 -120
rect 5575 -150 5625 -140
rect 5575 -170 5585 -150
rect 5605 -170 5625 -150
rect 5575 -175 5625 -170
rect 5680 -175 5700 -120
rect -20 -465 0 -300
rect -30 -485 0 -465
rect -240 -1150 -220 -485
rect 6440 -1085 6460 -80
rect 6925 -65 6975 -55
rect 6925 -85 6935 -65
rect 6955 -85 6975 -65
rect 6925 -90 6975 -85
rect 7030 -90 7050 45
rect 7995 -65 8045 -55
rect 7995 -85 8005 -65
rect 8025 -85 8045 -65
rect 7995 -90 8045 -85
rect 8100 -90 8120 45
rect 9065 -65 9115 -55
rect 9065 -85 9075 -65
rect 9095 -85 9115 -65
rect 9065 -90 9115 -85
rect 9170 -90 9190 45
rect 6680 -380 6700 -215
rect 6670 -400 6700 -380
rect 6440 -1105 6700 -1085
rect -240 -1160 -200 -1150
rect -240 -1180 -230 -1160
rect -210 -1170 -200 -1160
rect -210 -1180 0 -1170
rect -240 -1190 0 -1180
rect 7125 -1850 7165 -1840
rect 7125 -1870 7135 -1850
rect 7155 -1870 7165 -1850
rect 7125 -1880 7165 -1870
rect 7215 -1900 7235 -1840
rect 8195 -1850 8235 -1840
rect 8195 -1870 8205 -1850
rect 8225 -1870 8235 -1850
rect 8195 -1880 8235 -1870
rect 8285 -1900 8305 -1840
rect 9265 -1850 9305 -1840
rect 9265 -1870 9275 -1850
rect 9295 -1870 9305 -1850
rect 9265 -1880 9305 -1870
rect 9355 -1900 9375 -1840
rect 7215 -1920 9965 -1900
rect 425 -1935 465 -1925
rect 425 -1955 435 -1935
rect 455 -1955 465 -1935
rect 425 -1965 465 -1955
rect 515 -1985 535 -1925
rect 1495 -1935 1535 -1925
rect 1495 -1955 1505 -1935
rect 1525 -1955 1535 -1935
rect 1495 -1965 1535 -1955
rect 1585 -1985 1605 -1925
rect 2565 -1935 2605 -1925
rect 2565 -1955 2575 -1935
rect 2595 -1955 2605 -1935
rect 2565 -1965 2605 -1955
rect 2655 -1985 2675 -1925
rect 3635 -1935 3675 -1925
rect 3635 -1955 3645 -1935
rect 3665 -1955 3675 -1935
rect 3635 -1965 3675 -1955
rect 3725 -1985 3745 -1925
rect 4705 -1935 4745 -1925
rect 4705 -1955 4715 -1935
rect 4735 -1955 4745 -1935
rect 4705 -1965 4745 -1955
rect 4795 -1985 4815 -1925
rect 5775 -1935 5815 -1925
rect 5775 -1955 5785 -1935
rect 5805 -1955 5815 -1935
rect 5775 -1965 5815 -1955
rect 5865 -1985 5885 -1925
rect 9945 -1985 9965 -1920
rect 515 -2005 9965 -1985
rect -280 -2045 7490 -2025
rect -280 -3950 -260 -2045
rect 225 -2075 275 -2065
rect 225 -2095 235 -2075
rect 255 -2095 275 -2075
rect 225 -2100 275 -2095
rect 330 -2100 350 -2045
rect 1295 -2075 1345 -2065
rect 1295 -2095 1305 -2075
rect 1325 -2095 1345 -2075
rect 1295 -2100 1345 -2095
rect 1400 -2100 1420 -2045
rect 2365 -2075 2415 -2065
rect 2365 -2095 2375 -2075
rect 2395 -2095 2415 -2075
rect 2365 -2100 2415 -2095
rect 2470 -2100 2490 -2045
rect 3435 -2075 3485 -2065
rect 3435 -2095 3445 -2075
rect 3465 -2095 3485 -2075
rect 3435 -2100 3485 -2095
rect 3540 -2100 3560 -2045
rect 4505 -2075 4555 -2065
rect 4505 -2095 4515 -2075
rect 4535 -2095 4555 -2075
rect 4505 -2100 4555 -2095
rect 4610 -2100 4630 -2045
rect 5575 -2075 5625 -2065
rect 5575 -2095 5585 -2075
rect 5605 -2095 5625 -2075
rect 5575 -2100 5625 -2095
rect 5680 -2100 5700 -2045
rect 6645 -2075 6695 -2065
rect 6645 -2095 6655 -2075
rect 6675 -2095 6695 -2075
rect 6645 -2100 6695 -2095
rect 6750 -2100 6770 -2045
rect -20 -2390 0 -2225
rect -30 -2410 0 -2390
rect -240 -3075 -220 -2410
rect -240 -3085 -200 -3075
rect -240 -3105 -230 -3085
rect -210 -3095 -200 -3085
rect -210 -3105 0 -3095
rect -240 -3115 0 -3105
rect 425 -3860 465 -3850
rect 425 -3880 435 -3860
rect 455 -3880 465 -3860
rect 425 -3890 465 -3880
rect 515 -3910 535 -3850
rect 1495 -3860 1535 -3850
rect 1495 -3880 1505 -3860
rect 1525 -3880 1535 -3860
rect 1495 -3890 1535 -3880
rect 1585 -3910 1605 -3850
rect 2565 -3860 2605 -3850
rect 2565 -3880 2575 -3860
rect 2595 -3880 2605 -3860
rect 2565 -3890 2605 -3880
rect 2655 -3910 2675 -3850
rect 3635 -3860 3675 -3850
rect 3635 -3880 3645 -3860
rect 3665 -3880 3675 -3860
rect 3635 -3890 3675 -3880
rect 3725 -3910 3745 -3850
rect 4705 -3860 4745 -3850
rect 4705 -3880 4715 -3860
rect 4735 -3880 4745 -3860
rect 4705 -3890 4745 -3880
rect 4795 -3910 4815 -3850
rect 5775 -3860 5815 -3850
rect 5775 -3880 5785 -3860
rect 5805 -3880 5815 -3860
rect 5775 -3890 5815 -3880
rect 5865 -3910 5885 -3850
rect 6845 -3860 6885 -3850
rect 6845 -3880 6855 -3860
rect 6875 -3880 6885 -3860
rect 6845 -3890 6885 -3880
rect 6935 -3910 6955 -3850
rect 9945 -3910 9965 -2005
rect 515 -3930 9965 -3910
rect -280 -3970 7840 -3950
rect -280 -5875 -260 -3970
rect 225 -4000 275 -3990
rect 225 -4020 235 -4000
rect 255 -4020 275 -4000
rect 225 -4025 275 -4020
rect 330 -4025 350 -3970
rect 1295 -4000 1345 -3990
rect 1295 -4020 1305 -4000
rect 1325 -4020 1345 -4000
rect 1295 -4025 1345 -4020
rect 1400 -4025 1420 -3970
rect 2365 -4000 2415 -3990
rect 2365 -4020 2375 -4000
rect 2395 -4020 2415 -4000
rect 2365 -4025 2415 -4020
rect 2470 -4025 2490 -3970
rect 3435 -4000 3485 -3990
rect 3435 -4020 3445 -4000
rect 3465 -4020 3485 -4000
rect 3435 -4025 3485 -4020
rect 3540 -4025 3560 -3970
rect 4505 -4000 4555 -3990
rect 4505 -4020 4515 -4000
rect 4535 -4020 4555 -4000
rect 4505 -4025 4555 -4020
rect 4610 -4025 4630 -3970
rect 5575 -4000 5625 -3990
rect 5575 -4020 5585 -4000
rect 5605 -4020 5625 -4000
rect 5575 -4025 5625 -4020
rect 5680 -4025 5700 -3970
rect 6645 -4000 6695 -3990
rect 6645 -4020 6655 -4000
rect 6675 -4020 6695 -4000
rect 6645 -4025 6695 -4020
rect 6750 -4025 6770 -3970
rect 7715 -4000 7765 -3990
rect 7715 -4020 7725 -4000
rect 7745 -4020 7765 -4000
rect 7715 -4025 7765 -4020
rect 7820 -4025 7840 -3970
rect -20 -4315 0 -4150
rect -30 -4335 0 -4315
rect -240 -5000 -220 -4335
rect -240 -5010 -200 -5000
rect -240 -5030 -230 -5010
rect -210 -5020 -200 -5010
rect -210 -5030 0 -5020
rect -240 -5040 0 -5030
rect 425 -5785 465 -5775
rect 425 -5805 435 -5785
rect 455 -5805 465 -5785
rect 425 -5815 465 -5805
rect 515 -5835 535 -5775
rect 1495 -5785 1535 -5775
rect 1495 -5805 1505 -5785
rect 1525 -5805 1535 -5785
rect 1495 -5815 1535 -5805
rect 1585 -5835 1605 -5775
rect 2565 -5785 2605 -5775
rect 2565 -5805 2575 -5785
rect 2595 -5805 2605 -5785
rect 2565 -5815 2605 -5805
rect 2655 -5835 2675 -5775
rect 3635 -5785 3675 -5775
rect 3635 -5805 3645 -5785
rect 3665 -5805 3675 -5785
rect 3635 -5815 3675 -5805
rect 3725 -5835 3745 -5775
rect 4705 -5785 4745 -5775
rect 4705 -5805 4715 -5785
rect 4735 -5805 4745 -5785
rect 4705 -5815 4745 -5805
rect 4795 -5835 4815 -5775
rect 5775 -5785 5815 -5775
rect 5775 -5805 5785 -5785
rect 5805 -5805 5815 -5785
rect 5775 -5815 5815 -5805
rect 5865 -5835 5885 -5775
rect 6845 -5785 6885 -5775
rect 6845 -5805 6855 -5785
rect 6875 -5805 6885 -5785
rect 6845 -5815 6885 -5805
rect 6935 -5835 6955 -5775
rect 7915 -5785 7955 -5775
rect 7915 -5805 7925 -5785
rect 7945 -5805 7955 -5785
rect 7915 -5815 7955 -5805
rect 8005 -5835 8025 -5775
rect 9945 -5835 9965 -3930
rect 515 -5855 9965 -5835
rect -280 -5895 7490 -5875
rect -280 -7800 -260 -5895
rect 225 -5925 275 -5915
rect 225 -5945 235 -5925
rect 255 -5945 275 -5925
rect 225 -5950 275 -5945
rect 330 -5950 350 -5895
rect 1295 -5925 1345 -5915
rect 1295 -5945 1305 -5925
rect 1325 -5945 1345 -5925
rect 1295 -5950 1345 -5945
rect 1400 -5950 1420 -5895
rect 2365 -5925 2415 -5915
rect 2365 -5945 2375 -5925
rect 2395 -5945 2415 -5925
rect 2365 -5950 2415 -5945
rect 2470 -5950 2490 -5895
rect 3435 -5925 3485 -5915
rect 3435 -5945 3445 -5925
rect 3465 -5945 3485 -5925
rect 3435 -5950 3485 -5945
rect 3540 -5950 3560 -5895
rect 4505 -5925 4555 -5915
rect 4505 -5945 4515 -5925
rect 4535 -5945 4555 -5925
rect 4505 -5950 4555 -5945
rect 4610 -5950 4630 -5895
rect 5575 -5925 5625 -5915
rect 5575 -5945 5585 -5925
rect 5605 -5945 5625 -5925
rect 5575 -5950 5625 -5945
rect 5680 -5950 5700 -5895
rect 6645 -5925 6695 -5915
rect 6645 -5945 6655 -5925
rect 6675 -5945 6695 -5925
rect 6645 -5950 6695 -5945
rect 6750 -5950 6770 -5895
rect -20 -6240 0 -6075
rect -30 -6260 0 -6240
rect -240 -6925 -220 -6260
rect -240 -6935 -200 -6925
rect -240 -6955 -230 -6935
rect -210 -6945 -200 -6935
rect -210 -6955 0 -6945
rect -240 -6965 0 -6955
rect 425 -7710 465 -7700
rect 425 -7730 435 -7710
rect 455 -7730 465 -7710
rect 425 -7740 465 -7730
rect 515 -7760 535 -7700
rect 1495 -7710 1535 -7700
rect 1495 -7730 1505 -7710
rect 1525 -7730 1535 -7710
rect 1495 -7740 1535 -7730
rect 1585 -7760 1605 -7700
rect 2565 -7710 2605 -7700
rect 2565 -7730 2575 -7710
rect 2595 -7730 2605 -7710
rect 2565 -7740 2605 -7730
rect 2655 -7760 2675 -7700
rect 3635 -7710 3675 -7700
rect 3635 -7730 3645 -7710
rect 3665 -7730 3675 -7710
rect 3635 -7740 3675 -7730
rect 3725 -7760 3745 -7700
rect 4705 -7710 4745 -7700
rect 4705 -7730 4715 -7710
rect 4735 -7730 4745 -7710
rect 4705 -7740 4745 -7730
rect 4795 -7760 4815 -7700
rect 5775 -7710 5815 -7700
rect 5775 -7730 5785 -7710
rect 5805 -7730 5815 -7710
rect 5775 -7740 5815 -7730
rect 5865 -7760 5885 -7700
rect 6845 -7710 6885 -7700
rect 6845 -7730 6855 -7710
rect 6875 -7730 6885 -7710
rect 6845 -7740 6885 -7730
rect 6935 -7760 6955 -7700
rect 9945 -7760 9965 -5855
rect 515 -7780 9965 -7760
rect -280 -7820 9190 -7800
rect -340 -7850 -300 -7840
rect -340 -7870 -330 -7850
rect -310 -7870 -300 -7850
rect -340 -7880 -300 -7870
rect 225 -7850 275 -7840
rect 225 -7870 235 -7850
rect 255 -7870 275 -7850
rect 225 -7875 275 -7870
rect 330 -7875 350 -7820
rect 1295 -7850 1345 -7840
rect 1295 -7870 1305 -7850
rect 1325 -7870 1345 -7850
rect 1295 -7875 1345 -7870
rect 1400 -7875 1420 -7820
rect 2365 -7850 2415 -7840
rect 2365 -7870 2375 -7850
rect 2395 -7870 2415 -7850
rect 2365 -7875 2415 -7870
rect 2470 -7875 2490 -7820
rect 3435 -7850 3485 -7840
rect 3435 -7870 3445 -7850
rect 3465 -7870 3485 -7850
rect 3435 -7875 3485 -7870
rect 3540 -7875 3560 -7820
rect 4505 -7850 4555 -7840
rect 4505 -7870 4515 -7850
rect 4535 -7870 4555 -7850
rect 4505 -7875 4555 -7870
rect 4610 -7875 4630 -7820
rect 5575 -7850 5625 -7840
rect 5575 -7870 5585 -7850
rect 5605 -7870 5625 -7850
rect 5575 -7875 5625 -7870
rect 5680 -7875 5700 -7820
rect 6925 -7850 6975 -7840
rect 6925 -7870 6935 -7850
rect 6955 -7870 6975 -7850
rect 6925 -7875 6975 -7870
rect 7030 -7875 7050 -7820
rect 7995 -7850 8045 -7840
rect 7995 -7870 8005 -7850
rect 8025 -7870 8045 -7850
rect 7995 -7875 8045 -7870
rect 8100 -7875 8120 -7820
rect 9065 -7850 9115 -7840
rect 9065 -7870 9075 -7850
rect 9095 -7870 9115 -7850
rect 9065 -7875 9115 -7870
rect 9170 -7875 9190 -7820
rect -20 -8165 0 -8000
rect 6680 -8165 6700 -8000
rect -30 -8185 0 -8165
rect 6670 -8185 6700 -8165
rect -240 -8850 -220 -8185
rect -380 -8860 -340 -8850
rect -380 -8870 -370 -8860
rect -400 -8880 -370 -8870
rect -350 -8880 -340 -8860
rect -400 -8890 -340 -8880
rect -240 -8860 -200 -8850
rect -240 -8880 -230 -8860
rect -210 -8870 -200 -8860
rect 6460 -8870 6480 -8185
rect -210 -8880 0 -8870
rect -240 -8890 0 -8880
rect 6460 -8890 6700 -8870
rect 6460 -8975 6480 -8890
rect 6455 -9000 6480 -8975
rect 445 -9700 465 -9625
rect 425 -9710 465 -9700
rect 425 -9730 435 -9710
rect 455 -9730 465 -9710
rect 425 -9740 465 -9730
rect 515 -9765 535 -9625
rect 1515 -9700 1535 -9625
rect 1495 -9710 1535 -9700
rect 1495 -9730 1505 -9710
rect 1525 -9730 1535 -9710
rect 1495 -9740 1535 -9730
rect 1585 -9765 1605 -9625
rect 2585 -9700 2605 -9625
rect 2565 -9710 2605 -9700
rect 2565 -9730 2575 -9710
rect 2595 -9730 2605 -9710
rect 2565 -9740 2605 -9730
rect 2655 -9765 2675 -9625
rect 3655 -9700 3675 -9625
rect 3635 -9710 3675 -9700
rect 3635 -9730 3645 -9710
rect 3665 -9730 3675 -9710
rect 3635 -9740 3675 -9730
rect 3725 -9765 3745 -9625
rect 4725 -9700 4745 -9625
rect 4705 -9710 4745 -9700
rect 4705 -9730 4715 -9710
rect 4735 -9730 4745 -9710
rect 4705 -9740 4745 -9730
rect 4795 -9765 4815 -9625
rect 5795 -9700 5815 -9625
rect 5775 -9710 5815 -9700
rect 5775 -9730 5785 -9710
rect 5805 -9730 5815 -9710
rect 5775 -9740 5815 -9730
rect 5865 -9765 5885 -9625
rect 515 -9775 6430 -9765
rect 515 -9785 6400 -9775
rect 6390 -9795 6400 -9785
rect 6420 -9795 6430 -9775
rect 6390 -9805 6430 -9795
rect -380 -9815 -340 -9805
rect -380 -9825 -370 -9815
rect -400 -9835 -370 -9825
rect -350 -9835 -340 -9815
rect -400 -9845 -340 -9835
rect -240 -9815 -200 -9805
rect -240 -9835 -230 -9815
rect -210 -9825 -200 -9815
rect 6455 -9825 6475 -9000
rect 7125 -9635 7165 -9625
rect 7125 -9655 7135 -9635
rect 7155 -9655 7165 -9635
rect 7125 -9665 7165 -9655
rect 7215 -9685 7235 -9625
rect 8195 -9635 8235 -9625
rect 8195 -9655 8205 -9635
rect 8225 -9655 8235 -9635
rect 8195 -9665 8235 -9655
rect 8285 -9685 8305 -9625
rect 9265 -9635 9305 -9625
rect 9265 -9655 9275 -9635
rect 9295 -9655 9305 -9635
rect 9265 -9665 9305 -9655
rect 9355 -9685 9375 -9625
rect 9945 -9685 9965 -7780
rect 7215 -9705 9965 -9685
rect 9945 -9765 9965 -9705
rect 6695 -9775 9965 -9765
rect 6695 -9795 6705 -9775
rect 6725 -9785 9965 -9775
rect 6725 -9795 6735 -9785
rect 6695 -9805 6735 -9795
rect -210 -9835 6475 -9825
rect -240 -9845 6475 -9835
rect 9945 -9845 9965 -9785
rect 9985 -9795 10025 -9785
rect 9985 -9815 9995 -9795
rect 10015 -9805 10025 -9795
rect 10015 -9815 10045 -9805
rect 9985 -9825 10045 -9815
rect 9945 -9865 10045 -9845
<< metal1 >>
rect -290 -155 6460 -135
rect -290 -200 -270 -155
rect -290 -220 -240 -200
rect -290 -2125 -270 -220
rect -290 -2145 -235 -2125
rect -290 -4050 -270 -2145
rect -290 -4070 -235 -4050
rect -290 -5975 -270 -4070
rect -290 -5995 -235 -5975
rect -290 -7800 -270 -5995
rect -290 -7820 6490 -7800
rect -290 -7900 -270 -7820
rect 6460 -7900 6490 -7820
rect -290 -7920 -235 -7900
use dac_unit  dac_unit_0
timestamp 1702422646
transform 1 0 6825 0 1 -9645
box -125 20 945 1770
use dac_unit  dac_unit_1
timestamp 1702422646
transform 1 0 7895 0 1 -9645
box -125 20 945 1770
use dac_unit  dac_unit_2
timestamp 1702422646
transform 1 0 8965 0 1 -9645
box -125 20 945 1770
use dac_unit  dac_unit_3
timestamp 1702422646
transform 1 0 125 0 1 -1945
box -125 20 945 1770
use dac_unit  dac_unit_4
timestamp 1702422646
transform 1 0 1195 0 1 -1945
box -125 20 945 1770
use dac_unit  dac_unit_5
timestamp 1702422646
transform 1 0 2265 0 1 -1945
box -125 20 945 1770
use dac_unit  dac_unit_6
timestamp 1702422646
transform 1 0 3335 0 1 -1945
box -125 20 945 1770
use dac_unit  dac_unit_7
timestamp 1702422646
transform 1 0 4405 0 1 -1945
box -125 20 945 1770
use dac_unit  dac_unit_8
timestamp 1702422646
transform 1 0 5475 0 1 -1945
box -125 20 945 1770
use dac_unit  dac_unit_9
timestamp 1702422646
transform 1 0 125 0 1 -3870
box -125 20 945 1770
use dac_unit  dac_unit_10
timestamp 1702422646
transform 1 0 1195 0 1 -3870
box -125 20 945 1770
use dac_unit  dac_unit_11
timestamp 1702422646
transform 1 0 2265 0 1 -3870
box -125 20 945 1770
use dac_unit  dac_unit_12
timestamp 1702422646
transform 1 0 3335 0 1 -3870
box -125 20 945 1770
use dac_unit  dac_unit_13
timestamp 1702422646
transform 1 0 4405 0 1 -3870
box -125 20 945 1770
use dac_unit  dac_unit_14
timestamp 1702422646
transform 1 0 5475 0 1 -3870
box -125 20 945 1770
use dac_unit  dac_unit_15
timestamp 1702422646
transform 1 0 6545 0 1 -3870
box -125 20 945 1770
use dac_unit  dac_unit_16
timestamp 1702422646
transform 1 0 125 0 1 -5795
box -125 20 945 1770
use dac_unit  dac_unit_17
timestamp 1702422646
transform 1 0 1195 0 1 -5795
box -125 20 945 1770
use dac_unit  dac_unit_18
timestamp 1702422646
transform 1 0 2265 0 1 -5795
box -125 20 945 1770
use dac_unit  dac_unit_19
timestamp 1702422646
transform 1 0 3335 0 1 -5795
box -125 20 945 1770
use dac_unit  dac_unit_20
timestamp 1702422646
transform 1 0 4405 0 1 -5795
box -125 20 945 1770
use dac_unit  dac_unit_21
timestamp 1702422646
transform 1 0 5475 0 1 -5795
box -125 20 945 1770
use dac_unit  dac_unit_22
timestamp 1702422646
transform 1 0 6545 0 1 -5795
box -125 20 945 1770
use dac_unit  dac_unit_23
timestamp 1702422646
transform 1 0 7615 0 1 -5795
box -125 20 945 1770
use dac_unit  dac_unit_24
timestamp 1702422646
transform 1 0 125 0 1 -7720
box -125 20 945 1770
use dac_unit  dac_unit_25
timestamp 1702422646
transform 1 0 1195 0 1 -7720
box -125 20 945 1770
use dac_unit  dac_unit_26
timestamp 1702422646
transform 1 0 2265 0 1 -7720
box -125 20 945 1770
use dac_unit  dac_unit_27
timestamp 1702422646
transform 1 0 3335 0 1 -7720
box -125 20 945 1770
use dac_unit  dac_unit_28
timestamp 1702422646
transform 1 0 4405 0 1 -7720
box -125 20 945 1770
use dac_unit  dac_unit_29
timestamp 1702422646
transform 1 0 5475 0 1 -7720
box -125 20 945 1770
use dac_unit  dac_unit_30
timestamp 1702422646
transform 1 0 6545 0 1 -7720
box -125 20 945 1770
use dac_unit  dac_unit_31
timestamp 1702422646
transform 1 0 125 0 1 -9645
box -125 20 945 1770
use dac_unit  dac_unit_32
timestamp 1702422646
transform 1 0 1195 0 1 -9645
box -125 20 945 1770
use dac_unit  dac_unit_33
timestamp 1702422646
transform 1 0 2265 0 1 -9645
box -125 20 945 1770
use dac_unit  dac_unit_34
timestamp 1702422646
transform 1 0 3335 0 1 -9645
box -125 20 945 1770
use dac_unit  dac_unit_35
timestamp 1702422646
transform 1 0 4405 0 1 -9645
box -125 20 945 1770
use dac_unit  dac_unit_36
timestamp 1702422646
transform 1 0 5475 0 1 -9645
box -125 20 945 1770
use dac_unit  dac_unit_40
timestamp 1702422646
transform 1 0 6825 0 1 -1860
box -125 20 945 1770
use dac_unit  dac_unit_41
timestamp 1702422646
transform 1 0 7895 0 1 -1860
box -125 20 945 1770
use dac_unit  dac_unit_42
timestamp 1702422646
transform 1 0 8965 0 1 -1860
box -125 20 945 1770
use inverter  inverter_0
timestamp 1693780072
transform 1 0 6700 0 1 -8060
box -240 -145 -30 185
use inverter  inverter_1
timestamp 1693780072
transform 1 0 0 0 1 -360
box -240 -145 -30 185
use inverter  inverter_2
timestamp 1693780072
transform 1 0 0 0 1 -2285
box -240 -145 -30 185
use inverter  inverter_3
timestamp 1693780072
transform 1 0 0 0 1 -4210
box -240 -145 -30 185
use inverter  inverter_4
timestamp 1693780072
transform 1 0 0 0 1 -6135
box -240 -145 -30 185
use inverter  inverter_5
timestamp 1693780072
transform 1 0 0 0 1 -8060
box -240 -145 -30 185
use inverter  inverter_7
timestamp 1693780072
transform 1 0 6700 0 1 -275
box -240 -145 -30 185
<< labels >>
rlabel locali -400 -1180 -400 -1180 7 Vphi2
port 11 w
rlabel locali -400 -3105 -400 -3105 7 Vphi3
port 12 w
rlabel locali -400 -5030 -400 -5030 7 Vphi4
port 13 w
rlabel locali -400 -6955 -400 -6955 7 Vphi5
port 14 w
rlabel locali -400 -8880 -400 -8880 7 Vphi6
port 15 w
rlabel locali -400 -70 -400 -70 7 Vphi1
port 10 w
rlabel locali -400 55 -400 55 7 Vcp
port 8 w
rlabel locali -400 15 -400 15 7 Vbp
port 9 w
rlabel locali -400 -9835 -400 -9835 7 Vphi7
port 16 w
rlabel locali 10045 -9815 10045 -9815 3 Viout-
port 17 e
rlabel locali 10045 -9855 10045 -9855 3 Viout+
port 18 e
<< end >>
