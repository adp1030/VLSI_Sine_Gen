* NGSPICE file created from final.ext - technology: sky130A

.subckt v_gen VP VN Vb Vbp Vcp
X0 Vbp VP VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X1 Vcp Vb VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X2 a_740_1480# VP VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X3 a_1040_1370# a_1040_1370# a_940_1480# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X4 VN Vb a_740_1480# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X5 a_1040_1370# a_1040_1370# a_940_1480# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X6 VP a_1040_1370# a_940_1480# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X7 a_2330_1480# a_1040_1370# a_1040_1370# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X8 VP VP Vcp VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X9 VP VP Vbp VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X10 VN Vb a_2840_90# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X11 VN VN Vbp VN sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X12 a_1040_1370# a_1040_1370# a_2330_1480# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X13 a_1040_1370# a_1040_1370# a_2330_1480# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X14 VN Vb Vbp VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X15 a_2640_90# Vb a_2440_90# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X16 VN Vb Vb VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X17 a_2240_90# Vb a_1040_1370# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.65 ps=6.55 w=6 l=0.5
X18 a_1040_1370# Vb a_1830_90# VN sky130_fd_pr__nfet_01v8 ad=1.65 pd=6.55 as=1.5 ps=6.5 w=6 l=0.5
X19 a_1630_90# Vb a_1430_90# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X20 a_1230_90# Vb VN VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X21 VP Vbp Vbp VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X22 a_940_1480# a_740_1480# a_740_1480# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X23 a_940_1480# a_1040_1370# a_1040_1370# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X24 a_940_1480# a_1040_1370# a_1040_1370# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X25 Vcp Vcp a_2330_1480# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X26 Vbp Vbp VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X27 a_2330_1480# a_1040_1370# VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X28 Vbp Vb VN VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X29 a_2330_1480# a_1040_1370# a_1040_1370# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X30 Vb Vb VN VN sky130_fd_pr__nfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X31 a_2440_90# Vb a_2240_90# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X32 a_2840_90# Vb a_2640_90# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X33 Vbp VN VN VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X34 a_1830_90# Vb a_1630_90# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X35 a_1430_90# Vb a_1230_90# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
.ends

.subckt dac_unit Vbp Vcp Vphi Vphi_b Viup Viun VP
X0 a_3270_1770# Vcp a_2870_360# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X1 VP VP Viup VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X2 a_2870_360# Vcp a_2270_1770# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X3 Viun Vphi a_2870_360# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X4 a_2870_360# Vphi Viun VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X5 Viup VP VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X6 VP Vbp a_3270_1770# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=1.5 ps=6.5 w=6 l=0.5
X7 a_3270_1770# VP VP VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=3 ps=13 w=6 l=0.5
X8 VP VP a_2270_1770# VP sky130_fd_pr__pfet_01v8 ad=3 pd=13 as=3 ps=13 w=6 l=0.5
X9 a_2270_1770# Vbp VP VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=3 ps=13 w=6 l=0.5
X10 Viup Vphi_b a_2870_360# VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X11 a_2870_360# Vphi_b Viup VP sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
.ends

.subckt inverter A Y VP VN
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
.ends

.subckt dac Vcp VP Vphi1 VN Vphi7 Vphi5 Vphi2 Viout+ Vbp Viout- Vphi3 Vphi4 inverter_1/Y
+ Vphi6
Xdac_unit_4 Vbp Vcp Vphi2 inverter_2/Y Viout+ Viout- VP dac_unit
Xdac_unit_5 Vbp Vcp Vphi1 inverter_1/Y Viout+ Viout- VP dac_unit
Xdac_unit_6 Vbp Vcp Vphi5 inverter_5/Y Viout+ Viout- VP dac_unit
Xinverter_0 Vphi7 inverter_0/Y VP VN inverter
Xinverter_1 Vphi1 inverter_1/Y VP VN inverter
Xdac_unit_7 Vbp Vcp Vphi4 inverter_4/Y Viout+ Viout- VP dac_unit
Xinverter_2 Vphi2 inverter_2/Y VP VN inverter
Xdac_unit_8 Vbp Vcp Vphi4 inverter_4/Y Viout+ Viout- VP dac_unit
Xinverter_3 Vphi3 inverter_3/Y VP VN inverter
Xdac_unit_9 Vbp Vcp Vphi4 inverter_4/Y Viout+ Viout- VP dac_unit
Xinverter_4 Vphi4 inverter_4/Y VP VN inverter
Xinverter_5 Vphi5 inverter_5/Y VP VN inverter
Xinverter_6 Vphi6 inverter_6/Y VP VN inverter
Xdac_unit_40 Vbp Vcp Vphi1 inverter_1/Y Viout+ Viout- VP dac_unit
Xdac_unit_30 Vbp Vcp Vphi6 inverter_6/Y Viout+ Viout- VP dac_unit
Xdac_unit_20 Vbp Vcp Vphi5 inverter_5/Y Viout+ Viout- VP dac_unit
Xdac_unit_31 Vbp Vcp Vphi6 inverter_6/Y Viout+ Viout- VP dac_unit
Xdac_unit_21 Vbp Vcp Vphi3 inverter_3/Y Viout+ Viout- VP dac_unit
Xdac_unit_10 Vbp Vcp Vphi4 inverter_4/Y Viout+ Viout- VP dac_unit
Xdac_unit_32 Vbp Vcp Vphi6 inverter_6/Y Viout+ Viout- VP dac_unit
Xdac_unit_22 Vbp Vcp Vphi3 inverter_3/Y Viout+ Viout- VP dac_unit
Xdac_unit_11 Vbp Vcp Vphi4 inverter_4/Y Viout+ Viout- VP dac_unit
Xdac_unit_33 Vbp Vcp Vphi6 inverter_6/Y Viout+ Viout- VP dac_unit
Xdac_unit_23 Vbp Vcp Vphi3 inverter_3/Y Viout+ Viout- VP dac_unit
Xdac_unit_12 Vbp Vcp Vphi4 inverter_4/Y Viout+ Viout- VP dac_unit
Xdac_unit_34 Vbp Vcp Vphi6 inverter_6/Y Viout+ Viout- VP dac_unit
Xdac_unit_35 Vbp Vcp Vphi1 inverter_1/Y Viout+ Viout- VP dac_unit
Xdac_unit_13 Vbp Vcp Vphi2 inverter_2/Y Viout+ Viout- VP dac_unit
Xdac_unit_25 Vbp Vcp Vphi3 inverter_3/Y Viout+ Viout- VP dac_unit
Xdac_unit_24 Vbp Vcp Vphi3 inverter_3/Y Viout+ Viout- VP dac_unit
Xdac_unit_14 Vbp Vcp Vphi4 inverter_4/Y Viout+ Viout- VP dac_unit
Xdac_unit_36 Vbp Vcp Vphi7 inverter_0/Y Viout+ Viout- VP dac_unit
Xdac_unit_15 Vbp Vcp Vphi5 inverter_5/Y Viout+ Viout- VP dac_unit
Xdac_unit_37 Vbp Vcp Vphi7 inverter_0/Y Viout+ Viout- VP dac_unit
Xdac_unit_26 Vbp Vcp Vphi6 inverter_6/Y Viout+ Viout- VP dac_unit
Xdac_unit_27 Vbp Vcp Vphi3 inverter_3/Y Viout+ Viout- VP dac_unit
Xdac_unit_38 Vbp Vcp Vphi7 inverter_0/Y Viout+ Viout- VP dac_unit
Xdac_unit_16 Vbp Vcp Vphi5 inverter_5/Y Viout+ Viout- VP dac_unit
Xdac_unit_28 Vbp Vcp Vphi3 inverter_3/Y Viout+ Viout- VP dac_unit
Xdac_unit_17 Vbp Vcp Vphi5 inverter_5/Y Viout+ Viout- VP dac_unit
Xdac_unit_29 Vbp Vcp Vphi2 inverter_2/Y Viout+ Viout- VP dac_unit
Xdac_unit_18 Vbp Vcp Vphi5 inverter_5/Y Viout+ Viout- VP dac_unit
Xdac_unit_19 Vbp Vcp Vphi5 inverter_5/Y Viout+ Viout- VP dac_unit
Xdac_unit_0 Vbp Vcp Vphi4 inverter_4/Y Viout+ Viout- VP dac_unit
Xdac_unit_1 Vbp Vcp Vphi2 inverter_2/Y Viout+ Viout- VP dac_unit
Xdac_unit_3 Vbp Vcp Vphi2 inverter_2/Y Viout+ Viout- VP dac_unit
Xdac_unit_2 Vbp Vcp Vphi2 inverter_2/Y Viout+ Viout- VP dac_unit
.ends

.subckt filter VN Viout- Viout+
X0 Viout+ a_2360_6260# VN sky130_fd_pr__res_xhigh_po l=3.5
X1 VN a_2360_6260# VN sky130_fd_pr__res_xhigh_po l=3.5
X2 VN a_2360_1100# VN sky130_fd_pr__res_xhigh_po l=3.5
X3 a_1460_5820# a_1090_2450# sky130_fd_pr__cap_mim_m3_1 l=10 w=8
X4 Viout- a_2360_1100# VN sky130_fd_pr__res_xhigh_po l=3.5
X5 a_1460_5820# Vout+ VN sky130_fd_pr__res_xhigh_po l=3.5
X6 a_1090_2450# Viout- VN sky130_fd_pr__res_xhigh_po l=3.5
X7 a_1090_2450# Vout- VN sky130_fd_pr__res_xhigh_po l=3.5
X8 a_1460_5820# Viout+ VN sky130_fd_pr__res_xhigh_po l=3.5
X9 Vout+ Vout- sky130_fd_pr__cap_mim_m3_1 l=10 w=8
.ends

.subckt csrl_dff2 D DB Q QB CLK VP VN
X0 VP a_n950_630# a_n950_1180# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X1 a_n950_630# a_n950_1180# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X2 a_n950_630# CLK DB VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.75 ps=3.5 w=1 l=0.15
X3 QB CLK a_n950_630# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 VP a_n950_1180# a_n950_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X5 VN Q QB VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X6 a_n690_630# CLK VP VP sky130_fd_pr__pfet_01v8 ad=0.433 pd=3.03 as=0.5 ps=3.16 w=4 l=0.15
X7 a_n950_n280# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0.433 pd=3.03 as=2 ps=10.5 w=4 l=0.15
X8 a_n950_1180# a_n950_630# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X9 Q CLK a_n950_1180# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 VN QB Q VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X11 Q QB a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X12 QB Q a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X13 a_n950_1180# CLK D VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.75 ps=3.5 w=1 l=0.15
.ends

.subckt csrl_dff3 D DB Q QB CLK VP VN
X0 VP a_n950_630# a_n950_1180# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X1 a_n950_630# a_n950_1180# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X2 a_n950_630# CLK DB VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.75 ps=3.5 w=1 l=0.15
X3 QB CLK a_n950_630# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 VP a_n950_1180# a_n950_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X5 VN Q QB VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X6 a_n690_630# CLK VP VP sky130_fd_pr__pfet_01v8 ad=0.433 pd=3.03 as=0.5 ps=3.16 w=4 l=0.15
X7 a_n950_n280# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0.433 pd=3.03 as=2 ps=10.5 w=4 l=0.15
X8 a_n950_1180# a_n950_630# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X9 Q CLK a_n950_1180# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 VN QB Q VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X11 Q QB a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X12 QB Q a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X13 a_n950_1180# CLK D VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.75 ps=3.5 w=1 l=0.15
.ends

.subckt csrl_dff1 D DB Q QB CLK VP VN
X0 VP a_n950_630# a_n950_1180# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X1 a_n950_630# a_n950_1180# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X2 a_n950_630# CLK DB VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.55 ps=3.1 w=1 l=0.15
X3 QB CLK a_n950_630# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 VP a_n950_1180# a_n950_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3.16 as=0.25 ps=1.5 w=1 l=0.15
X5 VN Q QB VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X6 a_n690_630# CLK VP VP sky130_fd_pr__pfet_01v8 ad=0.433 pd=3.03 as=0.5 ps=3.16 w=4 l=0.15
X7 a_n950_n280# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0.433 pd=3.03 as=1.6 ps=9.7 w=4 l=0.15
X8 a_n950_1180# a_n950_630# a_n950_n280# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.433 ps=3.03 w=1 l=0.15
X9 Q CLK a_n950_1180# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X10 VN QB Q VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X11 Q QB a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X12 QB Q a_n690_630# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.433 ps=3.03 w=1 l=0.15
X13 a_n950_1180# CLK D VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.55 ps=3.1 w=1 l=0.15
.ends

.subckt register16 Vphi3 csrl_dff3_0/VP Vphi7 Vphi1 Vphi5 Vphi2 Vphi4 Vphi6 VSUBS
Xcsrl_dff2_10 csrl_dff2_9/Q csrl_dff2_9/QB csrl_dff2_11/D csrl_dff2_11/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_11 csrl_dff2_11/D csrl_dff2_11/DB csrl_dff2_12/D csrl_dff2_12/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_12 csrl_dff2_12/D csrl_dff2_12/DB csrl_dff2_13/D csrl_dff2_13/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_0 Vphi1 csrl_dff2_0/DB Vphi2 csrl_dff2_1/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_13 csrl_dff2_13/D csrl_dff2_13/DB csrl_dff3_0/D csrl_dff3_0/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_2 Vphi3 csrl_dff2_2/DB Vphi4 csrl_dff2_3/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_1 Vphi2 csrl_dff2_1/DB Vphi3 csrl_dff2_2/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_3 Vphi4 csrl_dff2_3/DB Vphi5 csrl_dff2_4/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_4 Vphi5 csrl_dff2_4/DB Vphi6 csrl_dff2_5/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_5 Vphi6 csrl_dff2_5/DB Vphi7 csrl_dff2_6/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_6 Vphi7 csrl_dff2_6/DB csrl_dff2_7/D csrl_dff2_7/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff2
Xcsrl_dff2_7 csrl_dff2_7/D csrl_dff2_7/DB csrl_dff2_8/D csrl_dff2_8/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_8 csrl_dff2_8/D csrl_dff2_8/DB csrl_dff2_9/D csrl_dff2_9/DB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff2_9 csrl_dff2_9/D csrl_dff2_9/DB csrl_dff2_9/Q csrl_dff2_9/QB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff2
Xcsrl_dff3_0 csrl_dff3_0/D csrl_dff3_0/DB csrl_dff3_0/Q csrl_dff3_0/QB csrl_dff3_0/CLK
+ csrl_dff3_0/VP VSUBS csrl_dff3
Xcsrl_dff1_0 csrl_dff3_0/Q csrl_dff3_0/QB Vphi1 csrl_dff2_0/DB csrl_dff3_0/CLK csrl_dff3_0/VP
+ VSUBS csrl_dff1
.ends


* Top level circuit final

Xv_gen_0 dac_0/VP VSUBS v_gen_0/Vb dac_0/Vbp dac_0/Vcp v_gen
Xdac_0 dac_0/Vcp dac_0/VP dac_0/Vphi1 VSUBS dac_0/Vphi7 dac_0/Vphi5 dac_0/Vphi2 dac_0/Viout+
+ dac_0/Vbp dac_0/Viout- dac_0/Vphi3 dac_0/Vphi4 dac_0/inverter_1/Y dac_0/Vphi6 dac
Xfilter_0 VSUBS dac_0/Viout- dac_0/Viout+ filter
Xregister16_0 dac_0/Vphi3 dac_0/VP dac_0/Vphi7 dac_0/Vphi1 dac_0/Vphi5 dac_0/Vphi2
+ dac_0/Vphi4 dac_0/Vphi6 VSUBS register16
.end

