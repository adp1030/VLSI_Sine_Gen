* NGSPICE file created from cap_test.ext - technology: sky130A


* Top level circuit cap_test

X0 top bot sky130_fd_pr__cap_mim_m3_1 l=10 w=8
X1 top bot sky130_fd_pr__cap_mim_m3_1 l=10 w=8
.end

