* NGSPICE file created from filter.ext - technology: sky130A

X0 a_n750_1380# Vout+ VN sky130_fd_pr__res_xhigh_po l=3.5
X1 a_n270_1030# VN VN sky130_fd_pr__res_xhigh_po l=3.5
X2 a_1640_1100# VN VN sky130_fd_pr__res_xhigh_po l=3.5
X3 a_2570_3400# Viout- VN sky130_fd_pr__res_xhigh_po l=3.5
X4 a_n270_1030# Viout+ VN sky130_fd_pr__res_xhigh_po l=3.5
X5 a_1640_1100# Viout- VN sky130_fd_pr__res_xhigh_po l=3.5
X6 Vout+ Vout- sky130_fd_pr__cap_mim_m3_1 l=10 w=8
X7 Vout- a_2570_3400# VN sky130_fd_pr__res_xhigh_po l=3.5
X8 a_n750_1380# Viout+ VN sky130_fd_pr__res_xhigh_po l=3.5
X9 a_n750_1380# a_2570_3400# sky130_fd_pr__cap_mim_m3_1 l=10 w=8
